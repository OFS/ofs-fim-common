// Copyright (C) 2023 Intel Corporation
// SPDX-License-Identifier: MIT

/**
 * Abstract: 
 * class 'pf_vf_mux_basic_env' is extended from uvm_env base class.  It implements
 * the build phase to construct the structural elements of this environment.
 *
 * pf_vf_mux_basic_env is the testbench environment, which constructs the AXI System
 * ENV in the build_phase method using the UVM factory service.  The AXI System
 * ENV  is the top level component provided by the AXI VIP. The AXI System ENV
 * in turn, instantiates constructs the AXI Master and Slave agents. 
 *
 * axi_basic env also constructs the virtual sequencer. This virtual sequencer
 * in the testbench environment obtains a handle to the reset interface using
 * the config db.  This allows reset sequences to be written for this virtual
 * sequencer.
 *
 * The simulation ends after all the objections are dropped.  This is done by
 * using objections provided by phase arguments.
 */
`ifndef GUARD_PF_VF_MUX_BASIC_ENV_SV
`define GUARD_PF_VF_MUX_BASIC_ENV_SV

`include "pf_vf_mux_scoreboard.sv"
`include "pf_vf_mux_virtual_sequencer.sv"

`define monitor_scoreboard_connection(PORT) \
  pf_vf_mux_system_env_H.master[0].monitor.item_observed_port.connect(pf_vf_mux_scbd_``PORT``.axi_port_rx);\
  pf_vf_mux_system_env_D.slave[``PORT``].monitor.item_observed_port.connect(pf_vf_mux_scbd_``PORT``.axi_port_tx);\

`define monitor_scoreboard_upstream_connection(PORT) \
  pf_vf_mux_system_env_H.slave[0].monitor.item_observed_port.connect(pf_vf_mux_scbd_``PORT``_up.axi_port_rx);\
  pf_vf_mux_system_env_D.master[``PORT``].monitor.item_observed_port.connect(pf_vf_mux_scbd_``PORT``_up.axi_port_tx);\

`define monitor_scoreboard_connection_N(VIP_PORT,RTL_PORT) \
  pf_vf_mux_system_env_H.master[0].monitor.item_observed_port.connect(pf_vf_mux_scbd_``RTL_PORT``.axi_port_rx);\
  pf_vf_mux_system_env_DN.slave[``VIP_PORT``].monitor.item_observed_port.connect(pf_vf_mux_scbd_``RTL_PORT``.axi_port_tx);\

`define monitor_scoreboard_upstream_connection_N(VIP_PORT,RTL_PORT) \
  pf_vf_mux_system_env_H.slave[0].monitor.item_observed_port.connect(pf_vf_mux_scbd_``RTL_PORT``_up.axi_port_rx);\
  pf_vf_mux_system_env_DN.master[``VIP_PORT``].monitor.item_observed_port.connect(pf_vf_mux_scbd_``RTL_PORT``_up.axi_port_tx);\

`define monitor_scoreboard_connection_TB4(VIP_NUM,RTL_PORT,VIP_PORT) \
  pf_vf_mux_system_env_H.master[0].monitor.item_observed_port.connect(pf_vf_mux_scbd_``RTL_PORT``.axi_port_rx);\
  pf_vf_mux_system_env_TB4_D``VIP_NUM``.slave[``VIP_PORT``].monitor.item_observed_port.connect(pf_vf_mux_scbd_``RTL_PORT``.axi_port_tx);\

`define monitor_scoreboard_upstream_connection_TB4(VIP_NUM,RTL_PORT,VIP_PORT) \
  pf_vf_mux_system_env_H.slave[0].monitor.item_observed_port.connect(pf_vf_mux_scbd_``RTL_PORT``_up.axi_port_rx);\
  pf_vf_mux_system_env_TB4_D``VIP_NUM``.master[``VIP_PORT``].monitor.item_observed_port.connect(pf_vf_mux_scbd_``RTL_PORT``_up.axi_port_tx);\


class pf_vf_mux_basic_env extends uvm_env;

  /** AXI System ENV */
  svt_axi_system_env   pf_vf_mux_system_env_H;
  svt_axi_system_env   pf_vf_mux_system_env_D;
  `ifndef TB_CONFIG_1
     `ifdef TB_CONFIG_4
       svt_axi_system_env   pf_vf_mux_system_env_TB4_D0;
       svt_axi_system_env   pf_vf_mux_system_env_TB4_D1;
       svt_axi_system_env   pf_vf_mux_system_env_TB4_D2;
       svt_axi_system_env   pf_vf_mux_system_env_TB4_D3;
     `else  
       svt_axi_system_env   pf_vf_mux_system_env_DN;
     `endif  
  `endif

  pf_vf_mux_scoreboard  pf_vf_mux_scbd_0;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_3;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_4;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_5;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_6;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_7;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_8;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_9;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_10;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_11;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_12;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_13;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_14;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_15;
  `ifdef TB_CONFIG_2
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_16;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_17;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_18;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_19;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_20;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_21;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_22;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_23;
  `elsif TB_CONFIG_3
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_16;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_17;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_18;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_19;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_20;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_21;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_22;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_23;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_24;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_25;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_26;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_27;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_28;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_29;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_30;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_31;
  `elsif TB_CONFIG_4
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_16;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_17;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_18;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_19;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_20;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_21;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_22;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_23;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_24;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_25;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_26;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_27;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_28;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_29;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_30;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_31;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_32;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_33;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_34;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_35;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_36;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_37;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_38;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_39;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_40;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_41;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_42;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_43;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_44;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_45;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_46;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_47;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_48;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_49;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_50;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_51;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_52;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_53;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_54;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_55;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_56;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_57;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_58;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_59;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_60;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_61;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_62;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_63;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_64;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_65;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_66;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_67;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_68;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_69;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_70;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_71;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_72;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_73;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_74;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_75;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_76;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_77;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_78;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_79;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_80;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_81;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_82;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_83;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_84;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_85;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_86;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_87;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_88;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_89;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_90;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_91;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_92;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_93;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_94;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_95;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_96;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_97;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_98;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_99;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_100;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_101;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_102;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_103;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_104;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_105;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_106;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_107;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_108;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_109;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_110;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_111;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_112;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_113;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_114;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_115;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_116;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_117;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_118;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_119;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_120;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_121;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_122;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_123;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_124;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_125;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_126;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_127;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_128;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_129;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_130;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_131;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_132;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_133;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_134;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_135;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_136;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_137;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_138;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_139;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_140;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_141;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_142;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_143;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_144;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_145;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_146;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_147;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_148;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_149;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_150;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_151;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_152;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_153;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_154;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_155;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_156;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_157;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_158;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_159;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_160;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_161;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_162;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_163;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_164;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_165;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_166;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_167;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_168;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_169;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_170;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_171;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_172;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_173;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_174;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_175;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_176;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_177;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_178;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_179;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_180;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_181;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_182;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_183;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_184;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_185;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_186;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_187;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_188;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_189;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_190;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_191;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_192;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_193;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_194;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_195;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_196;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_197;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_198;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_199;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_200;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_201;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_202;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_203;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_204;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_205;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_206;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_207;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_208;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_209;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_210;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_211;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_212;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_213;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_214;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_215;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_216;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_217;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_218;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_219;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_220;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_221;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_222;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_223;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_224;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_225;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_226;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_227;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_228;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_229;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_230;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_231;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_232;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_233;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_234;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_235;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_236;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_237;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_238;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_239;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_240;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_241;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_242;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_243;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_244;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_245;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_246;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_247;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_248;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_249;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_250;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_251;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_252;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_253;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_254;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_255;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_256;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_257;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_258;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_259;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_260;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_261;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_262;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_263;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_264;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_265;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_266;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_267;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_268;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_269;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_270;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_271;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_272;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_273;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_274;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_275;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_276;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_277;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_278;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_279;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_280;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_281;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_282;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_283;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_284;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_285;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_286;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_287;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_288;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_289;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_290;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_291;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_292;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_293;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_294;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_295;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_296;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_297;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_298;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_299;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_300;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_301;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_302;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_303;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_304;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_305;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_306;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_307;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_308;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_309;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_310;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_311;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_312;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_313;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_314;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_315;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_316;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_317;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_318;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_319;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_320;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_321;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_322;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_323;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_324;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_325;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_326;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_327;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_328;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_329;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_330;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_331;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_332;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_333;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_334;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_335;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_336;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_337;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_338;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_339;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_340;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_341;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_342;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_343;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_344;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_345;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_346;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_347;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_348;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_349;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_350;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_351;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_352;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_353;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_354;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_355;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_356;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_357;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_358;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_359;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_360;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_361;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_362;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_363;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_364;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_365;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_366;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_367;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_368;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_369;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_370;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_371;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_372;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_373;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_374;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_375;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_376;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_377;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_378;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_379;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_380;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_381;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_382;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_383;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_384;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_385;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_386;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_387;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_388;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_389;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_390;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_391;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_392;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_393;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_394;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_395;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_396;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_397;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_398;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_399;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_400;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_401;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_402;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_403;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_404;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_405;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_406;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_407;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_408;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_409;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_410;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_411;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_412;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_413;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_414;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_415;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_416;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_417;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_418;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_419;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_420;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_421;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_422;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_423;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_424;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_425;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_426;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_427;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_428;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_429;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_430;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_431;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_432;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_433;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_434;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_435;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_436;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_437;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_438;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_439;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_440;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_441;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_442;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_443;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_444;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_445;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_446;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_447;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_448;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_449;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_450;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_451;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_452;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_453;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_454;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_455;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_456;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_457;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_458;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_459;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_460;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_461;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_462;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_463;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_464;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_465;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_466;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_467;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_468;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_469;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_470;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_471;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_472;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_473;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_474;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_475;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_476;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_477;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_478;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_479;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_480;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_481;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_482;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_483;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_484;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_485;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_486;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_487;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_488;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_489;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_490;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_491;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_492;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_493;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_494;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_495;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_496;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_497;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_498;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_499;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_500;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_501;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_502;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_503;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_504;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_505;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_506;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_507;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_508;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_509;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_510;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_511;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_512;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_513;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_514;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_515;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_516;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_517;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_518;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_519;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_520;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_521;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_522;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_523;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_524;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_525;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_526;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_527;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_528;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_529;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_530;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_531;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_532;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_533;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_534;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_535;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_536;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_537;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_538;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_539;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_540;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_541;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_542;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_543;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_544;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_545;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_546;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_547;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_548;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_549;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_550;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_551;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_552;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_553;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_554;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_555;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_556;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_557;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_558;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_559;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_560;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_561;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_562;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_563;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_564;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_565;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_566;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_567;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_568;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_569;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_570;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_571;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_572;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_573;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_574;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_575;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_576;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_577;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_578;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_579;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_580;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_581;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_582;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_583;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_584;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_585;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_586;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_587;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_588;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_589;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_590;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_591;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_592;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_593;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_594;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_595;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_596;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_597;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_598;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_599;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_600;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_601;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_602;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_603;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_604;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_605;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_606;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_607;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_608;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_609;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_610;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_611;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_612;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_613;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_614;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_615;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_616;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_617;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_618;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_619;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_620;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_621;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_622;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_623;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_624;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_625;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_626;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_627;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_628;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_629;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_630;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_631;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_632;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_633;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_634;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_635;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_636;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_637;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_638;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_639;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_640;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_641;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_642;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_643;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_644;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_645;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_646;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_647;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_648;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_649;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_650;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_651;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_652;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_653;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_654;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_655;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_656;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_657;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_658;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_659;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_660;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_661;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_662;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_663;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_664;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_665;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_666;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_667;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_668;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_669;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_670;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_671;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_672;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_673;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_674;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_675;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_676;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_677;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_678;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_679;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_680;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_681;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_682;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_683;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_684;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_685;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_686;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_687;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_688;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_689;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_690;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_691;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_692;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_693;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_694;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_695;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_696;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_697;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_698;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_699;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_700;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_701;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_702;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_703;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_704;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_705;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_706;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_707;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_708;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_709;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_710;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_711;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_712;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_713;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_714;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_715;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_716;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_717;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_718;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_719;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_720;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_721;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_722;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_723;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_724;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_725;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_726;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_727;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_728;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_729;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_730;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_731;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_732;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_733;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_734;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_735;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_736;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_737;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_738;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_739;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_740;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_741;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_742;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_743;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_744;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_745;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_746;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_747;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_748;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_749;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_750;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_751;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_752;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_753;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_754;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_755;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_756;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_757;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_758;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_759;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_760;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_761;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_762;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_763;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_764;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_765;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_766;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_767;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_768;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_769;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_770;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_771;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_772;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_773;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_774;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_775;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_776;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_777;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_778;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_779;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_780;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_781;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_782;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_783;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_784;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_785;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_786;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_787;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_788;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_789;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_790;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_791;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_792;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_793;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_794;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_795;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_796;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_797;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_798;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_799;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_800;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_801;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_802;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_803;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_804;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_805;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_806;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_807;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_808;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_809;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_810;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_811;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_812;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_813;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_814;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_815;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_816;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_817;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_818;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_819;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_820;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_821;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_822;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_823;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_824;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_825;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_826;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_827;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_828;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_829;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_830;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_831;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_832;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_833;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_834;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_835;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_836;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_837;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_838;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_839;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_840;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_841;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_842;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_843;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_844;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_845;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_846;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_847;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_848;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_849;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_850;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_851;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_852;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_853;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_854;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_855;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_856;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_857;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_858;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_859;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_860;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_861;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_862;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_863;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_864;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_865;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_866;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_867;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_868;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_869;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_870;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_871;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_872;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_873;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_874;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_875;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_876;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_877;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_878;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_879;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_880;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_881;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_882;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_883;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_884;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_885;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_886;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_887;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_888;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_889;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_890;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_891;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_892;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_893;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_894;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_895;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_896;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_897;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_898;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_899;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_900;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_901;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_902;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_903;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_904;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_905;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_906;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_907;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_908;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_909;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_910;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_911;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_912;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_913;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_914;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_915;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_916;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_917;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_918;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_919;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_920;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_921;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_922;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_923;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_924;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_925;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_926;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_927;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_928;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_929;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_930;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_931;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_932;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_933;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_934;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_935;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_936;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_937;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_938;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_939;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_940;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_941;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_942;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_943;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_944;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_945;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_946;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_947;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_948;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_949;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_950;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_951;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_952;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_953;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_954;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_955;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_956;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_957;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_958;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_959;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_960;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_961;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_962;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_963;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_964;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_965;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_966;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_967;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_968;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_969;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_970;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_971;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_972;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_973;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_974;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_975;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_976;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_977;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_978;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_979;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_980;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_981;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_982;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_983;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_984;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_985;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_986;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_987;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_988;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_989;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_990;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_991;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_992;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_993;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_994;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_995;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_996;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_997;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_998;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_999;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1000;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1001;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1002;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1003;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1004;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1005;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1006;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1007;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1008;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1009;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1010;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1011;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1012;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1013;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1014;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1015;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1016;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1017;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1018;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1019;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1020;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1021;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1022;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1023;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1024;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1025;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1026;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1027;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1028;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1029;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1030;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1031;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1032;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1033;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1034;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1035;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1036;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1037;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1038;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1039;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1040;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1041;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1042;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1043;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1044;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1045;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1046;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1047;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1048;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1049;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1050;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1051;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1052;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1053;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1054;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1055;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1056;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1057;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1058;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1059;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1060;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1061;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1062;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1063;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1064;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1065;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1066;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1067;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1068;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1069;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1070;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1071;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1072;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1073;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1074;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1075;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1076;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1077;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1078;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1079;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1080;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1081;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1082;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1083;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1084;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1085;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1086;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1087;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1088;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1089;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1090;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1091;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1092;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1093;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1094;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1095;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1096;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1097;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1098;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1099;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1100;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1101;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1102;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1103;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1104;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1105;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1106;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1107;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1108;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1109;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1110;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1111;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1112;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1113;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1114;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1115;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1116;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1117;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1118;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1119;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1120;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1121;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1122;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1123;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1124;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1125;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1126;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1127;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1128;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1129;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1130;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1131;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1132;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1133;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1134;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1135;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1136;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1137;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1138;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1139;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1140;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1141;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1142;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1143;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1144;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1145;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1146;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1147;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1148;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1149;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1150;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1151;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1152;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1153;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1154;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1155;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1156;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1157;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1158;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1159;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1160;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1161;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1162;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1163;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1164;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1165;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1166;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1167;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1168;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1169;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1170;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1171;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1172;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1173;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1174;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1175;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1176;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1177;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1178;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1179;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1180;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1181;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1182;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1183;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1184;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1185;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1186;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1187;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1188;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1189;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1190;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1191;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1192;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1193;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1194;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1195;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1196;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1197;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1198;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1199;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1200;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1201;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1202;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1203;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1204;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1205;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1206;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1207;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1208;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1209;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1210;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1211;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1212;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1213;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1214;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1215;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1216;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1217;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1218;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1219;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1220;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1221;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1222;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1223;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1224;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1225;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1226;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1227;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1228;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1229;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1230;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1231;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1232;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1233;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1234;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1235;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1236;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1237;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1238;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1239;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1240;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1241;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1242;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1243;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1244;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1245;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1246;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1247;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1248;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1249;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1250;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1251;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1252;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1253;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1254;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1255;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1256;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1257;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1258;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1259;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1260;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1261;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1262;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1263;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1264;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1265;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1266;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1267;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1268;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1269;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1270;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1271;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1272;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1273;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1274;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1275;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1276;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1277;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1278;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1279;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1280;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1281;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1282;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1283;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1284;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1285;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1286;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1287;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1288;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1289;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1290;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1291;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1292;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1293;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1294;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1295;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1296;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1297;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1298;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1299;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1300;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1301;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1302;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1303;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1304;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1305;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1306;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1307;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1308;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1309;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1310;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1311;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1312;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1313;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1314;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1315;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1316;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1317;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1318;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1319;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1320;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1321;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1322;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1323;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1324;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1325;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1326;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1327;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1328;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1329;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1330;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1331;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1332;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1333;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1334;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1335;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1336;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1337;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1338;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1339;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1340;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1341;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1342;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1343;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1344;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1345;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1346;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1347;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1348;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1349;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1350;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1351;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1352;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1353;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1354;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1355;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1356;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1357;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1358;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1359;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1360;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1361;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1362;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1363;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1364;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1365;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1366;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1367;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1368;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1369;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1370;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1371;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1372;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1373;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1374;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1375;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1376;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1377;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1378;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1379;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1380;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1381;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1382;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1383;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1384;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1385;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1386;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1387;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1388;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1389;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1390;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1391;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1392;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1393;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1394;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1395;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1396;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1397;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1398;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1399;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1400;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1401;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1402;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1403;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1404;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1405;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1406;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1407;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1408;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1409;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1410;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1411;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1412;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1413;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1414;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1415;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1416;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1417;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1418;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1419;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1420;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1421;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1422;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1423;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1424;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1425;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1426;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1427;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1428;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1429;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1430;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1431;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1432;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1433;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1434;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1435;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1436;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1437;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1438;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1439;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1440;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1441;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1442;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1443;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1444;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1445;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1446;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1447;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1448;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1449;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1450;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1451;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1452;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1453;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1454;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1455;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1456;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1457;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1458;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1459;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1460;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1461;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1462;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1463;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1464;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1465;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1466;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1467;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1468;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1469;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1470;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1471;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1472;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1473;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1474;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1475;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1476;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1477;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1478;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1479;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1480;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1481;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1482;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1483;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1484;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1485;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1486;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1487;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1488;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1489;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1490;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1491;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1492;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1493;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1494;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1495;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1496;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1497;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1498;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1499;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1500;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1501;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1502;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1503;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1504;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1505;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1506;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1507;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1508;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1509;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1510;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1511;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1512;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1513;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1514;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1515;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1516;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1517;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1518;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1519;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1520;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1521;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1522;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1523;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1524;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1525;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1526;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1527;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1528;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1529;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1530;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1531;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1532;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1533;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1534;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1535;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1536;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1537;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1538;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1539;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1540;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1541;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1542;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1543;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1544;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1545;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1546;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1547;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1548;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1549;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1550;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1551;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1552;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1553;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1554;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1555;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1556;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1557;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1558;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1559;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1560;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1561;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1562;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1563;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1564;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1565;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1566;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1567;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1568;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1569;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1570;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1571;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1572;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1573;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1574;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1575;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1576;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1577;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1578;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1579;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1580;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1581;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1582;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1583;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1584;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1585;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1586;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1587;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1588;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1589;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1590;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1591;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1592;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1593;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1594;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1595;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1596;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1597;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1598;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1599;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1600;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1601;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1602;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1603;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1604;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1605;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1606;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1607;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1608;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1609;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1610;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1611;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1612;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1613;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1614;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1615;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1616;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1617;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1618;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1619;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1620;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1621;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1622;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1623;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1624;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1625;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1626;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1627;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1628;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1629;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1630;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1631;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1632;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1633;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1634;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1635;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1636;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1637;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1638;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1639;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1640;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1641;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1642;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1643;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1644;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1645;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1646;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1647;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1648;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1649;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1650;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1651;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1652;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1653;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1654;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1655;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1656;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1657;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1658;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1659;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1660;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1661;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1662;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1663;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1664;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1665;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1666;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1667;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1668;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1669;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1670;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1671;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1672;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1673;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1674;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1675;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1676;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1677;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1678;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1679;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1680;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1681;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1682;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1683;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1684;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1685;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1686;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1687;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1688;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1689;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1690;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1691;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1692;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1693;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1694;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1695;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1696;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1697;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1698;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1699;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1700;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1701;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1702;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1703;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1704;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1705;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1706;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1707;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1708;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1709;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1710;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1711;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1712;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1713;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1714;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1715;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1716;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1717;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1718;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1719;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1720;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1721;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1722;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1723;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1724;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1725;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1726;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1727;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1728;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1729;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1730;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1731;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1732;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1733;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1734;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1735;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1736;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1737;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1738;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1739;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1740;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1741;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1742;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1743;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1744;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1745;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1746;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1747;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1748;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1749;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1750;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1751;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1752;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1753;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1754;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1755;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1756;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1757;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1758;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1759;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1760;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1761;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1762;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1763;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1764;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1765;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1766;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1767;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1768;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1769;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1770;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1771;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1772;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1773;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1774;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1775;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1776;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1777;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1778;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1779;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1780;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1781;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1782;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1783;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1784;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1785;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1786;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1787;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1788;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1789;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1790;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1791;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1792;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1793;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1794;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1795;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1796;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1797;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1798;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1799;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1800;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1801;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1802;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1803;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1804;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1805;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1806;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1807;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1808;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1809;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1810;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1811;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1812;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1813;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1814;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1815;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1816;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1817;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1818;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1819;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1820;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1821;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1822;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1823;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1824;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1825;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1826;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1827;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1828;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1829;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1830;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1831;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1832;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1833;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1834;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1835;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1836;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1837;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1838;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1839;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1840;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1841;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1842;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1843;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1844;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1845;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1846;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1847;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1848;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1849;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1850;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1851;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1852;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1853;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1854;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1855;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1856;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1857;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1858;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1859;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1860;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1861;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1862;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1863;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1864;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1865;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1866;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1867;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1868;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1869;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1870;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1871;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1872;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1873;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1874;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1875;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1876;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1877;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1878;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1879;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1880;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1881;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1882;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1883;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1884;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1885;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1886;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1887;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1888;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1889;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1890;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1891;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1892;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1893;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1894;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1895;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1896;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1897;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1898;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1899;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1900;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1901;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1902;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1903;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1904;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1905;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1906;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1907;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1908;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1909;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1910;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1911;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1912;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1913;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1914;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1915;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1916;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1917;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1918;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1919;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1920;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1921;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1922;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1923;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1924;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1925;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1926;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1927;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1928;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1929;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1930;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1931;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1932;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1933;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1934;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1935;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1936;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1937;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1938;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1939;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1940;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1941;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1942;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1943;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1944;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1945;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1946;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1947;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1948;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1949;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1950;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1951;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1952;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1953;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1954;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1955;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1956;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1957;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1958;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1959;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1960;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1961;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1962;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1963;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1964;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1965;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1966;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1967;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1968;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1969;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1970;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1971;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1972;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1973;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1974;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1975;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1976;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1977;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1978;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1979;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1980;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1981;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1982;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1983;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1984;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1985;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1986;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1987;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1988;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1989;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1990;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1991;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1992;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1993;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1994;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1995;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1996;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1997;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1998;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1999;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2000;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2001;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2002;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2003;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2004;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2005;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2006;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2007;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2008;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2009;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2010;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2011;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2012;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2013;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2014;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2015;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2016;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2017;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2018;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2019;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2020;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2021;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2022;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2023;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2024;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2025;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2026;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2027;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2028;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2029;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2030;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2031;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2032;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2033;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2034;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2035;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2036;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2037;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2038;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2039;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2040;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2041;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2042;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2043;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2044;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2045;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2046;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2047;
  `endif
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_0_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_3_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_4_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_5_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_6_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_7_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_8_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_9_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_10_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_11_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_12_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_13_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_14_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_15_up;
  `ifdef TB_CONFIG_2
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_16_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_17_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_18_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_19_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_20_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_21_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_22_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_23_up;
  `elsif TB_CONFIG_3
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_16_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_17_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_18_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_19_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_20_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_21_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_22_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_23_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_24_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_25_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_26_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_27_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_28_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_29_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_30_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_31_up;
  `elsif TB_CONFIG_4
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_16_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_17_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_18_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_19_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_20_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_21_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_22_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_23_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_24_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_25_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_26_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_27_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_28_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_29_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_30_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_31_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_32_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_33_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_34_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_35_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_36_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_37_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_38_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_39_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_40_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_41_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_42_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_43_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_44_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_45_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_46_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_47_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_48_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_49_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_50_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_51_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_52_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_53_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_54_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_55_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_56_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_57_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_58_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_59_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_60_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_61_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_62_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_63_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_64_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_65_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_66_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_67_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_68_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_69_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_70_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_71_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_72_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_73_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_74_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_75_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_76_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_77_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_78_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_79_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_80_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_81_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_82_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_83_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_84_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_85_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_86_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_87_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_88_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_89_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_90_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_91_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_92_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_93_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_94_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_95_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_96_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_97_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_98_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_99_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_100_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_101_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_102_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_103_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_104_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_105_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_106_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_107_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_108_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_109_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_110_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_111_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_112_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_113_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_114_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_115_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_116_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_117_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_118_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_119_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_120_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_121_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_122_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_123_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_124_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_125_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_126_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_127_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_128_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_129_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_130_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_131_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_132_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_133_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_134_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_135_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_136_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_137_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_138_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_139_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_140_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_141_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_142_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_143_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_144_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_145_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_146_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_147_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_148_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_149_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_150_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_151_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_152_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_153_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_154_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_155_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_156_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_157_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_158_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_159_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_160_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_161_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_162_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_163_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_164_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_165_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_166_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_167_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_168_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_169_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_170_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_171_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_172_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_173_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_174_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_175_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_176_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_177_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_178_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_179_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_180_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_181_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_182_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_183_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_184_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_185_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_186_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_187_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_188_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_189_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_190_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_191_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_192_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_193_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_194_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_195_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_196_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_197_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_198_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_199_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_200_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_201_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_202_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_203_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_204_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_205_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_206_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_207_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_208_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_209_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_210_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_211_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_212_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_213_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_214_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_215_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_216_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_217_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_218_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_219_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_220_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_221_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_222_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_223_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_224_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_225_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_226_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_227_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_228_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_229_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_230_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_231_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_232_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_233_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_234_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_235_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_236_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_237_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_238_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_239_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_240_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_241_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_242_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_243_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_244_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_245_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_246_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_247_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_248_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_249_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_250_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_251_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_252_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_253_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_254_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_255_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_256_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_257_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_258_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_259_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_260_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_261_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_262_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_263_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_264_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_265_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_266_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_267_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_268_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_269_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_270_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_271_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_272_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_273_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_274_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_275_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_276_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_277_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_278_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_279_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_280_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_281_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_282_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_283_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_284_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_285_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_286_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_287_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_288_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_289_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_290_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_291_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_292_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_293_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_294_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_295_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_296_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_297_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_298_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_299_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_300_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_301_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_302_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_303_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_304_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_305_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_306_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_307_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_308_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_309_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_310_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_311_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_312_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_313_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_314_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_315_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_316_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_317_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_318_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_319_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_320_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_321_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_322_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_323_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_324_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_325_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_326_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_327_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_328_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_329_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_330_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_331_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_332_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_333_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_334_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_335_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_336_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_337_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_338_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_339_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_340_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_341_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_342_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_343_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_344_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_345_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_346_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_347_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_348_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_349_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_350_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_351_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_352_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_353_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_354_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_355_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_356_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_357_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_358_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_359_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_360_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_361_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_362_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_363_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_364_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_365_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_366_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_367_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_368_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_369_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_370_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_371_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_372_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_373_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_374_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_375_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_376_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_377_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_378_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_379_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_380_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_381_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_382_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_383_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_384_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_385_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_386_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_387_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_388_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_389_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_390_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_391_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_392_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_393_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_394_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_395_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_396_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_397_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_398_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_399_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_400_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_401_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_402_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_403_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_404_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_405_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_406_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_407_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_408_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_409_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_410_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_411_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_412_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_413_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_414_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_415_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_416_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_417_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_418_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_419_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_420_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_421_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_422_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_423_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_424_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_425_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_426_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_427_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_428_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_429_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_430_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_431_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_432_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_433_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_434_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_435_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_436_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_437_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_438_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_439_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_440_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_441_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_442_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_443_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_444_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_445_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_446_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_447_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_448_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_449_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_450_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_451_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_452_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_453_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_454_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_455_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_456_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_457_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_458_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_459_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_460_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_461_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_462_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_463_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_464_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_465_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_466_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_467_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_468_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_469_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_470_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_471_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_472_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_473_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_474_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_475_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_476_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_477_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_478_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_479_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_480_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_481_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_482_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_483_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_484_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_485_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_486_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_487_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_488_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_489_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_490_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_491_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_492_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_493_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_494_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_495_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_496_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_497_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_498_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_499_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_500_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_501_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_502_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_503_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_504_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_505_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_506_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_507_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_508_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_509_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_510_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_511_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_512_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_513_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_514_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_515_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_516_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_517_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_518_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_519_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_520_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_521_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_522_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_523_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_524_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_525_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_526_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_527_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_528_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_529_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_530_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_531_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_532_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_533_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_534_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_535_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_536_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_537_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_538_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_539_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_540_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_541_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_542_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_543_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_544_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_545_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_546_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_547_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_548_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_549_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_550_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_551_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_552_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_553_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_554_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_555_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_556_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_557_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_558_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_559_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_560_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_561_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_562_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_563_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_564_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_565_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_566_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_567_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_568_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_569_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_570_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_571_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_572_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_573_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_574_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_575_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_576_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_577_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_578_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_579_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_580_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_581_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_582_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_583_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_584_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_585_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_586_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_587_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_588_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_589_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_590_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_591_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_592_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_593_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_594_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_595_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_596_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_597_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_598_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_599_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_600_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_601_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_602_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_603_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_604_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_605_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_606_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_607_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_608_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_609_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_610_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_611_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_612_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_613_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_614_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_615_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_616_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_617_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_618_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_619_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_620_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_621_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_622_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_623_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_624_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_625_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_626_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_627_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_628_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_629_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_630_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_631_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_632_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_633_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_634_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_635_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_636_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_637_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_638_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_639_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_640_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_641_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_642_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_643_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_644_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_645_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_646_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_647_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_648_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_649_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_650_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_651_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_652_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_653_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_654_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_655_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_656_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_657_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_658_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_659_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_660_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_661_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_662_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_663_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_664_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_665_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_666_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_667_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_668_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_669_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_670_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_671_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_672_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_673_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_674_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_675_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_676_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_677_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_678_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_679_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_680_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_681_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_682_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_683_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_684_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_685_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_686_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_687_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_688_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_689_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_690_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_691_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_692_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_693_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_694_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_695_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_696_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_697_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_698_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_699_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_700_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_701_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_702_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_703_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_704_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_705_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_706_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_707_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_708_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_709_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_710_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_711_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_712_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_713_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_714_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_715_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_716_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_717_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_718_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_719_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_720_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_721_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_722_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_723_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_724_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_725_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_726_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_727_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_728_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_729_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_730_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_731_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_732_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_733_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_734_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_735_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_736_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_737_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_738_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_739_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_740_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_741_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_742_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_743_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_744_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_745_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_746_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_747_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_748_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_749_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_750_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_751_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_752_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_753_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_754_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_755_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_756_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_757_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_758_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_759_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_760_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_761_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_762_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_763_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_764_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_765_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_766_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_767_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_768_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_769_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_770_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_771_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_772_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_773_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_774_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_775_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_776_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_777_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_778_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_779_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_780_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_781_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_782_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_783_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_784_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_785_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_786_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_787_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_788_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_789_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_790_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_791_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_792_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_793_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_794_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_795_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_796_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_797_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_798_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_799_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_800_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_801_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_802_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_803_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_804_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_805_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_806_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_807_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_808_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_809_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_810_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_811_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_812_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_813_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_814_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_815_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_816_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_817_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_818_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_819_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_820_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_821_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_822_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_823_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_824_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_825_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_826_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_827_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_828_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_829_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_830_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_831_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_832_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_833_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_834_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_835_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_836_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_837_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_838_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_839_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_840_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_841_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_842_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_843_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_844_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_845_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_846_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_847_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_848_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_849_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_850_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_851_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_852_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_853_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_854_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_855_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_856_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_857_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_858_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_859_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_860_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_861_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_862_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_863_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_864_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_865_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_866_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_867_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_868_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_869_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_870_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_871_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_872_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_873_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_874_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_875_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_876_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_877_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_878_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_879_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_880_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_881_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_882_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_883_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_884_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_885_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_886_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_887_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_888_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_889_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_890_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_891_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_892_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_893_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_894_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_895_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_896_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_897_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_898_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_899_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_900_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_901_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_902_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_903_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_904_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_905_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_906_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_907_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_908_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_909_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_910_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_911_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_912_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_913_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_914_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_915_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_916_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_917_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_918_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_919_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_920_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_921_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_922_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_923_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_924_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_925_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_926_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_927_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_928_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_929_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_930_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_931_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_932_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_933_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_934_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_935_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_936_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_937_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_938_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_939_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_940_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_941_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_942_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_943_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_944_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_945_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_946_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_947_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_948_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_949_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_950_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_951_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_952_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_953_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_954_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_955_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_956_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_957_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_958_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_959_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_960_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_961_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_962_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_963_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_964_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_965_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_966_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_967_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_968_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_969_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_970_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_971_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_972_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_973_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_974_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_975_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_976_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_977_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_978_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_979_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_980_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_981_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_982_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_983_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_984_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_985_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_986_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_987_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_988_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_989_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_990_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_991_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_992_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_993_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_994_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_995_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_996_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_997_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_998_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_999_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1000_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1001_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1002_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1003_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1004_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1005_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1006_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1007_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1008_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1009_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1010_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1011_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1012_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1013_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1014_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1015_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1016_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1017_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1018_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1019_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1020_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1021_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1022_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1023_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1024_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1025_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1026_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1027_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1028_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1029_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1030_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1031_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1032_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1033_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1034_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1035_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1036_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1037_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1038_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1039_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1040_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1041_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1042_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1043_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1044_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1045_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1046_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1047_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1048_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1049_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1050_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1051_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1052_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1053_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1054_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1055_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1056_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1057_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1058_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1059_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1060_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1061_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1062_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1063_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1064_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1065_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1066_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1067_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1068_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1069_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1070_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1071_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1072_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1073_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1074_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1075_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1076_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1077_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1078_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1079_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1080_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1081_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1082_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1083_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1084_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1085_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1086_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1087_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1088_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1089_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1090_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1091_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1092_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1093_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1094_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1095_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1096_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1097_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1098_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1099_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1100_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1101_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1102_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1103_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1104_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1105_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1106_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1107_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1108_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1109_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1110_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1111_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1112_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1113_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1114_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1115_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1116_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1117_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1118_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1119_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1120_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1121_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1122_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1123_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1124_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1125_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1126_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1127_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1128_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1129_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1130_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1131_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1132_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1133_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1134_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1135_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1136_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1137_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1138_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1139_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1140_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1141_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1142_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1143_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1144_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1145_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1146_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1147_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1148_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1149_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1150_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1151_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1152_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1153_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1154_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1155_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1156_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1157_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1158_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1159_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1160_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1161_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1162_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1163_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1164_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1165_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1166_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1167_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1168_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1169_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1170_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1171_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1172_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1173_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1174_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1175_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1176_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1177_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1178_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1179_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1180_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1181_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1182_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1183_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1184_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1185_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1186_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1187_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1188_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1189_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1190_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1191_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1192_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1193_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1194_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1195_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1196_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1197_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1198_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1199_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1200_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1201_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1202_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1203_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1204_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1205_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1206_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1207_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1208_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1209_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1210_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1211_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1212_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1213_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1214_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1215_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1216_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1217_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1218_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1219_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1220_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1221_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1222_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1223_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1224_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1225_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1226_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1227_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1228_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1229_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1230_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1231_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1232_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1233_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1234_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1235_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1236_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1237_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1238_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1239_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1240_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1241_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1242_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1243_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1244_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1245_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1246_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1247_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1248_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1249_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1250_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1251_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1252_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1253_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1254_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1255_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1256_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1257_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1258_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1259_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1260_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1261_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1262_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1263_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1264_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1265_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1266_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1267_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1268_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1269_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1270_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1271_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1272_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1273_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1274_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1275_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1276_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1277_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1278_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1279_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1280_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1281_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1282_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1283_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1284_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1285_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1286_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1287_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1288_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1289_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1290_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1291_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1292_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1293_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1294_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1295_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1296_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1297_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1298_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1299_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1300_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1301_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1302_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1303_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1304_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1305_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1306_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1307_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1308_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1309_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1310_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1311_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1312_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1313_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1314_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1315_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1316_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1317_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1318_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1319_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1320_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1321_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1322_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1323_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1324_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1325_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1326_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1327_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1328_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1329_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1330_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1331_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1332_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1333_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1334_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1335_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1336_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1337_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1338_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1339_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1340_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1341_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1342_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1343_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1344_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1345_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1346_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1347_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1348_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1349_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1350_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1351_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1352_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1353_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1354_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1355_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1356_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1357_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1358_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1359_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1360_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1361_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1362_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1363_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1364_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1365_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1366_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1367_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1368_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1369_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1370_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1371_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1372_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1373_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1374_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1375_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1376_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1377_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1378_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1379_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1380_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1381_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1382_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1383_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1384_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1385_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1386_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1387_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1388_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1389_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1390_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1391_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1392_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1393_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1394_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1395_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1396_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1397_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1398_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1399_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1400_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1401_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1402_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1403_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1404_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1405_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1406_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1407_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1408_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1409_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1410_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1411_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1412_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1413_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1414_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1415_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1416_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1417_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1418_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1419_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1420_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1421_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1422_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1423_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1424_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1425_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1426_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1427_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1428_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1429_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1430_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1431_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1432_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1433_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1434_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1435_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1436_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1437_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1438_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1439_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1440_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1441_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1442_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1443_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1444_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1445_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1446_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1447_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1448_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1449_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1450_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1451_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1452_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1453_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1454_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1455_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1456_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1457_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1458_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1459_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1460_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1461_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1462_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1463_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1464_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1465_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1466_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1467_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1468_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1469_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1470_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1471_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1472_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1473_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1474_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1475_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1476_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1477_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1478_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1479_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1480_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1481_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1482_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1483_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1484_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1485_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1486_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1487_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1488_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1489_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1490_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1491_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1492_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1493_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1494_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1495_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1496_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1497_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1498_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1499_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1500_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1501_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1502_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1503_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1504_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1505_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1506_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1507_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1508_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1509_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1510_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1511_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1512_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1513_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1514_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1515_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1516_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1517_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1518_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1519_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1520_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1521_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1522_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1523_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1524_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1525_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1526_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1527_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1528_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1529_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1530_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1531_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1532_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1533_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1534_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1535_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1536_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1537_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1538_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1539_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1540_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1541_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1542_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1543_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1544_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1545_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1546_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1547_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1548_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1549_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1550_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1551_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1552_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1553_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1554_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1555_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1556_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1557_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1558_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1559_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1560_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1561_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1562_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1563_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1564_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1565_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1566_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1567_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1568_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1569_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1570_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1571_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1572_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1573_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1574_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1575_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1576_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1577_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1578_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1579_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1580_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1581_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1582_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1583_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1584_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1585_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1586_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1587_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1588_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1589_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1590_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1591_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1592_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1593_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1594_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1595_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1596_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1597_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1598_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1599_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1600_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1601_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1602_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1603_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1604_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1605_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1606_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1607_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1608_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1609_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1610_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1611_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1612_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1613_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1614_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1615_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1616_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1617_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1618_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1619_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1620_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1621_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1622_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1623_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1624_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1625_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1626_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1627_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1628_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1629_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1630_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1631_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1632_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1633_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1634_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1635_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1636_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1637_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1638_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1639_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1640_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1641_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1642_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1643_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1644_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1645_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1646_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1647_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1648_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1649_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1650_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1651_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1652_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1653_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1654_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1655_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1656_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1657_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1658_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1659_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1660_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1661_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1662_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1663_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1664_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1665_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1666_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1667_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1668_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1669_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1670_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1671_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1672_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1673_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1674_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1675_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1676_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1677_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1678_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1679_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1680_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1681_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1682_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1683_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1684_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1685_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1686_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1687_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1688_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1689_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1690_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1691_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1692_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1693_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1694_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1695_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1696_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1697_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1698_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1699_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1700_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1701_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1702_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1703_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1704_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1705_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1706_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1707_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1708_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1709_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1710_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1711_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1712_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1713_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1714_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1715_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1716_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1717_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1718_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1719_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1720_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1721_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1722_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1723_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1724_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1725_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1726_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1727_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1728_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1729_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1730_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1731_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1732_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1733_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1734_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1735_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1736_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1737_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1738_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1739_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1740_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1741_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1742_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1743_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1744_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1745_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1746_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1747_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1748_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1749_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1750_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1751_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1752_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1753_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1754_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1755_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1756_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1757_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1758_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1759_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1760_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1761_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1762_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1763_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1764_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1765_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1766_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1767_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1768_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1769_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1770_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1771_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1772_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1773_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1774_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1775_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1776_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1777_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1778_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1779_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1780_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1781_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1782_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1783_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1784_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1785_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1786_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1787_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1788_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1789_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1790_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1791_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1792_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1793_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1794_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1795_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1796_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1797_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1798_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1799_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1800_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1801_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1802_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1803_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1804_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1805_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1806_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1807_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1808_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1809_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1810_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1811_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1812_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1813_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1814_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1815_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1816_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1817_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1818_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1819_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1820_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1821_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1822_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1823_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1824_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1825_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1826_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1827_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1828_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1829_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1830_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1831_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1832_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1833_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1834_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1835_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1836_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1837_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1838_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1839_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1840_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1841_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1842_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1843_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1844_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1845_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1846_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1847_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1848_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1849_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1850_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1851_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1852_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1853_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1854_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1855_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1856_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1857_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1858_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1859_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1860_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1861_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1862_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1863_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1864_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1865_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1866_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1867_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1868_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1869_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1870_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1871_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1872_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1873_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1874_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1875_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1876_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1877_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1878_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1879_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1880_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1881_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1882_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1883_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1884_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1885_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1886_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1887_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1888_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1889_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1890_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1891_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1892_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1893_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1894_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1895_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1896_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1897_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1898_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1899_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1900_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1901_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1902_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1903_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1904_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1905_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1906_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1907_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1908_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1909_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1910_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1911_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1912_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1913_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1914_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1915_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1916_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1917_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1918_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1919_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1920_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1921_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1922_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1923_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1924_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1925_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1926_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1927_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1928_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1929_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1930_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1931_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1932_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1933_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1934_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1935_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1936_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1937_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1938_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1939_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1940_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1941_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1942_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1943_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1944_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1945_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1946_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1947_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1948_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1949_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1950_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1951_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1952_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1953_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1954_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1955_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1956_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1957_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1958_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1959_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1960_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1961_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1962_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1963_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1964_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1965_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1966_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1967_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1968_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1969_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1970_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1971_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1972_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1973_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1974_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1975_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1976_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1977_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1978_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1979_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1980_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1981_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1982_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1983_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1984_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1985_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1986_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1987_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1988_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1989_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1990_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1991_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1992_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1993_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1994_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1995_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1996_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1997_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1998_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_1999_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2000_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2001_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2002_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2003_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2004_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2005_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2006_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2007_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2008_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2009_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2010_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2011_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2012_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2013_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2014_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2015_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2016_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2017_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2018_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2019_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2020_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2021_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2022_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2023_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2024_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2025_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2026_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2027_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2028_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2029_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2030_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2031_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2032_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2033_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2034_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2035_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2036_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2037_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2038_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2039_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2040_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2041_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2042_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2043_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2044_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2045_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2046_up;
  pf_vf_mux_scoreboard  pf_vf_mux_scbd_2047_up;
  `endif


  /** Virtual Sequencer */
  pf_vf_mux_virtual_sequencer sequencer;

  /** AXI System Configuration */
  svt_axi_system_configuration cfg_H;
  svt_axi_system_configuration cfg_D;
  `ifndef TB_CONFIG_1
    `ifdef TB_CONFIG_4
       svt_axi_system_configuration cfg_TB4_D0;
       svt_axi_system_configuration cfg_TB4_D1;
       svt_axi_system_configuration cfg_TB4_D2;
       svt_axi_system_configuration cfg_TB4_D3;
    `else
       svt_axi_system_configuration cfg_DN;
     `endif
  `endif

  /** UVM Component Utility macro */
  `uvm_component_utils(pf_vf_mux_basic_env)

  /** Class Constructor */
  function new (string name="pf_vf_mux_basic_env", uvm_component parent=null);
    super.new (name, parent);
  endfunction

  /** Build the AXI System ENV */
  virtual function void build_phase(uvm_phase phase);
    `uvm_info("build_phase", "Entered...",UVM_LOW)

    super.build_phase(phase);

      cfg_H = svt_axi_system_configuration::type_id::create("cfg_H");
      cfg_D = svt_axi_system_configuration::type_id::create("cfg_D");
      AXIS_HOST_CFG();
      AXIS_DEVICE_CFG();
      `ifndef TB_CONFIG_1
         `ifdef TB_CONFIG_4
           cfg_TB4_D0 = svt_axi_system_configuration::type_id::create("cfg_TB4_D0");
           cfg_TB4_D1 = svt_axi_system_configuration::type_id::create("cfg_TB4_D1");
           cfg_TB4_D2 = svt_axi_system_configuration::type_id::create("cfg_TB4_D2");
           cfg_TB4_D3 = svt_axi_system_configuration::type_id::create("cfg_TB4_D3");
			     AXIS_DEVICE_TB4_CFG();
         `else
            cfg_DN = svt_axi_system_configuration::type_id::create("cfg_DN");
            AXIS_DEVICE_CFG_N();
          `endif  
       `endif
      /** Apply the configuration to the System ENV */
      uvm_config_db#(svt_axi_system_configuration)::set(this, "pf_vf_mux_system_env_H", "cfg", cfg_H);
      uvm_config_db#(svt_axi_system_configuration)::set(this, "pf_vf_mux_system_env_D", "cfg", cfg_D);
      `ifndef TB_CONFIG_1
         `ifdef TB_CONFIG_4
            uvm_config_db#(svt_axi_system_configuration)::set(this, "pf_vf_mux_system_env_TB4_D0", "cfg", cfg_TB4_D0);
      uvm_config_db#(svt_axi_system_configuration)::set(this, "pf_vf_mux_system_env_TB4_D1", "cfg", cfg_TB4_D1);
      uvm_config_db#(svt_axi_system_configuration)::set(this, "pf_vf_mux_system_env_TB4_D2", "cfg", cfg_TB4_D2);
      uvm_config_db#(svt_axi_system_configuration)::set(this, "pf_vf_mux_system_env_TB4_D3", "cfg", cfg_TB4_D3);
         `else
            uvm_config_db#(svt_axi_system_configuration)::set(this, "pf_vf_mux_system_env_DN", "cfg", cfg_DN);
           `endif 
      `endif
      // end

    /** Construct the system agent */
    pf_vf_mux_system_env_H = svt_axi_system_env::type_id::create("pf_vf_mux_system_env_H", this);
    pf_vf_mux_system_env_D = svt_axi_system_env::type_id::create("pf_vf_mux_system_env_D", this);
      `ifndef TB_CONFIG_1
         `ifdef TB_CONFIG_4
            pf_vf_mux_system_env_TB4_D0 = svt_axi_system_env::type_id::create("pf_vf_mux_system_env_TB4_D0", this);
            pf_vf_mux_system_env_TB4_D1 = svt_axi_system_env::type_id::create("pf_vf_mux_system_env_TB4_D1", this);
            pf_vf_mux_system_env_TB4_D2 = svt_axi_system_env::type_id::create("pf_vf_mux_system_env_TB4_D2", this);
            pf_vf_mux_system_env_TB4_D3 = svt_axi_system_env::type_id::create("pf_vf_mux_system_env_TB4_D3", this);
         `else
            pf_vf_mux_system_env_DN = svt_axi_system_env::type_id::create("pf_vf_mux_system_env_DN", this);
      `endif
    `endif
    pf_vf_mux_scbd_0 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_0", this);
    pf_vf_mux_scbd_1 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1", this);
    pf_vf_mux_scbd_2 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2", this);
    pf_vf_mux_scbd_3 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_3", this);
    pf_vf_mux_scbd_4 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_4", this);
    pf_vf_mux_scbd_5 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_5", this);
    pf_vf_mux_scbd_6 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_6", this);
    pf_vf_mux_scbd_7 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_7", this);
    pf_vf_mux_scbd_8 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_8", this);
    pf_vf_mux_scbd_9 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_9", this);
    pf_vf_mux_scbd_10 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_10", this);
    pf_vf_mux_scbd_11 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_11", this);
    pf_vf_mux_scbd_12 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_12", this);
    pf_vf_mux_scbd_13 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_13", this);
    pf_vf_mux_scbd_14 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_14", this);
    pf_vf_mux_scbd_15 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_15", this);
    `ifdef TB_CONFIG_2
    pf_vf_mux_scbd_16 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_16", this);
    pf_vf_mux_scbd_17 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_17", this);
    pf_vf_mux_scbd_18 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_18", this);
    pf_vf_mux_scbd_19 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_19", this);
    pf_vf_mux_scbd_20 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_20", this);
    pf_vf_mux_scbd_21 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_21", this);
    pf_vf_mux_scbd_22 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_22", this);
    pf_vf_mux_scbd_23 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_23", this);
    `elsif TB_CONFIG_3
    pf_vf_mux_scbd_16 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_16", this);
    pf_vf_mux_scbd_17 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_17", this);
    pf_vf_mux_scbd_18 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_18", this);
    pf_vf_mux_scbd_19 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_19", this);
    pf_vf_mux_scbd_20 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_20", this);
    pf_vf_mux_scbd_21 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_21", this);
    pf_vf_mux_scbd_22 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_22", this);
    pf_vf_mux_scbd_23 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_23", this);
    pf_vf_mux_scbd_24 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_24", this);
    pf_vf_mux_scbd_25 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_25", this);
    pf_vf_mux_scbd_26 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_26", this);
    pf_vf_mux_scbd_27 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_27", this);
    pf_vf_mux_scbd_28 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_28", this);
    pf_vf_mux_scbd_29 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_29", this);
    pf_vf_mux_scbd_30 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_30", this);
    pf_vf_mux_scbd_31 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_31", this);
    `elsif TB_CONFIG_4
    pf_vf_mux_scbd_16 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_16", this);
    pf_vf_mux_scbd_17 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_17", this);
    pf_vf_mux_scbd_18 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_18", this);
    pf_vf_mux_scbd_19 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_19", this);
    pf_vf_mux_scbd_20 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_20", this);
    pf_vf_mux_scbd_21 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_21", this);
    pf_vf_mux_scbd_22 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_22", this);
    pf_vf_mux_scbd_23 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_23", this);
    pf_vf_mux_scbd_24 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_24", this);
    pf_vf_mux_scbd_25 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_25", this);
    pf_vf_mux_scbd_26 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_26", this);
    pf_vf_mux_scbd_27 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_27", this);
    pf_vf_mux_scbd_28 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_28", this);
    pf_vf_mux_scbd_29 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_29", this);
    pf_vf_mux_scbd_30 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_30", this);
    pf_vf_mux_scbd_31 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_31", this);
    pf_vf_mux_scbd_32 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_32", this);
    pf_vf_mux_scbd_33 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_33", this);
    pf_vf_mux_scbd_34 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_34", this);
    pf_vf_mux_scbd_35 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_35", this);
    pf_vf_mux_scbd_36 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_36", this);
    pf_vf_mux_scbd_37 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_37", this);
    pf_vf_mux_scbd_38 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_38", this);
    pf_vf_mux_scbd_39 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_39", this);
    pf_vf_mux_scbd_40 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_40", this);
    pf_vf_mux_scbd_41 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_41", this);
    pf_vf_mux_scbd_42 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_42", this);
    pf_vf_mux_scbd_43 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_43", this);
    pf_vf_mux_scbd_44 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_44", this);
    pf_vf_mux_scbd_45 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_45", this);
    pf_vf_mux_scbd_46 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_46", this);
    pf_vf_mux_scbd_47 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_47", this);
    pf_vf_mux_scbd_48 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_48", this);
    pf_vf_mux_scbd_49 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_49", this);
    pf_vf_mux_scbd_50 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_50", this);
    pf_vf_mux_scbd_51 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_51", this);
    pf_vf_mux_scbd_52 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_52", this);
    pf_vf_mux_scbd_53 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_53", this);
    pf_vf_mux_scbd_54 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_54", this);
    pf_vf_mux_scbd_55 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_55", this);
    pf_vf_mux_scbd_56 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_56", this);
    pf_vf_mux_scbd_57 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_57", this);
    pf_vf_mux_scbd_58 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_58", this);
    pf_vf_mux_scbd_59 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_59", this);
    pf_vf_mux_scbd_60 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_60", this);
    pf_vf_mux_scbd_61 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_61", this);
    pf_vf_mux_scbd_62 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_62", this);
    pf_vf_mux_scbd_63 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_63", this);
    pf_vf_mux_scbd_64 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_64", this);
    pf_vf_mux_scbd_65 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_65", this);
    pf_vf_mux_scbd_66 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_66", this);
    pf_vf_mux_scbd_67 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_67", this);
    pf_vf_mux_scbd_68 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_68", this);
    pf_vf_mux_scbd_69 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_69", this);
    pf_vf_mux_scbd_70 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_70", this);
    pf_vf_mux_scbd_71 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_71", this);
    pf_vf_mux_scbd_72 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_72", this);
    pf_vf_mux_scbd_73 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_73", this);
    pf_vf_mux_scbd_74 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_74", this);
    pf_vf_mux_scbd_75 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_75", this);
    pf_vf_mux_scbd_76 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_76", this);
    pf_vf_mux_scbd_77 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_77", this);
    pf_vf_mux_scbd_78 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_78", this);
    pf_vf_mux_scbd_79 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_79", this);
    pf_vf_mux_scbd_80 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_80", this);
    pf_vf_mux_scbd_81 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_81", this);
    pf_vf_mux_scbd_82 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_82", this);
    pf_vf_mux_scbd_83 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_83", this);
    pf_vf_mux_scbd_84 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_84", this);
    pf_vf_mux_scbd_85 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_85", this);
    pf_vf_mux_scbd_86 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_86", this);
    pf_vf_mux_scbd_87 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_87", this);
    pf_vf_mux_scbd_88 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_88", this);
    pf_vf_mux_scbd_89 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_89", this);
    pf_vf_mux_scbd_90 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_90", this);
    pf_vf_mux_scbd_91 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_91", this);
    pf_vf_mux_scbd_92 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_92", this);
    pf_vf_mux_scbd_93 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_93", this);
    pf_vf_mux_scbd_94 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_94", this);
    pf_vf_mux_scbd_95 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_95", this);
    pf_vf_mux_scbd_96 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_96", this);
    pf_vf_mux_scbd_97 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_97", this);
    pf_vf_mux_scbd_98 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_98", this);
    pf_vf_mux_scbd_99 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_99", this);
    pf_vf_mux_scbd_100 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_100", this);
    pf_vf_mux_scbd_101 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_101", this);
    pf_vf_mux_scbd_102 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_102", this);
    pf_vf_mux_scbd_103 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_103", this);
    pf_vf_mux_scbd_104 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_104", this);
    pf_vf_mux_scbd_105 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_105", this);
    pf_vf_mux_scbd_106 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_106", this);
    pf_vf_mux_scbd_107 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_107", this);
    pf_vf_mux_scbd_108 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_108", this);
    pf_vf_mux_scbd_109 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_109", this);
    pf_vf_mux_scbd_110 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_110", this);
    pf_vf_mux_scbd_111 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_111", this);
    pf_vf_mux_scbd_112 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_112", this);
    pf_vf_mux_scbd_113 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_113", this);
    pf_vf_mux_scbd_114 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_114", this);
    pf_vf_mux_scbd_115 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_115", this);
    pf_vf_mux_scbd_116 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_116", this);
    pf_vf_mux_scbd_117 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_117", this);
    pf_vf_mux_scbd_118 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_118", this);
    pf_vf_mux_scbd_119 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_119", this);
    pf_vf_mux_scbd_120 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_120", this);
    pf_vf_mux_scbd_121 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_121", this);
    pf_vf_mux_scbd_122 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_122", this);
    pf_vf_mux_scbd_123 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_123", this);
    pf_vf_mux_scbd_124 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_124", this);
    pf_vf_mux_scbd_125 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_125", this);
    pf_vf_mux_scbd_126 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_126", this);
    pf_vf_mux_scbd_127 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_127", this);
    pf_vf_mux_scbd_128 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_128", this);
    pf_vf_mux_scbd_129 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_129", this);
    pf_vf_mux_scbd_130 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_130", this);
    pf_vf_mux_scbd_131 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_131", this);
    pf_vf_mux_scbd_132 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_132", this);
    pf_vf_mux_scbd_133 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_133", this);
    pf_vf_mux_scbd_134 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_134", this);
    pf_vf_mux_scbd_135 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_135", this);
    pf_vf_mux_scbd_136 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_136", this);
    pf_vf_mux_scbd_137 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_137", this);
    pf_vf_mux_scbd_138 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_138", this);
    pf_vf_mux_scbd_139 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_139", this);
    pf_vf_mux_scbd_140 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_140", this);
    pf_vf_mux_scbd_141 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_141", this);
    pf_vf_mux_scbd_142 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_142", this);
    pf_vf_mux_scbd_143 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_143", this);
    pf_vf_mux_scbd_144 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_144", this);
    pf_vf_mux_scbd_145 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_145", this);
    pf_vf_mux_scbd_146 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_146", this);
    pf_vf_mux_scbd_147 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_147", this);
    pf_vf_mux_scbd_148 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_148", this);
    pf_vf_mux_scbd_149 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_149", this);
    pf_vf_mux_scbd_150 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_150", this);
    pf_vf_mux_scbd_151 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_151", this);
    pf_vf_mux_scbd_152 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_152", this);
    pf_vf_mux_scbd_153 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_153", this);
    pf_vf_mux_scbd_154 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_154", this);
    pf_vf_mux_scbd_155 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_155", this);
    pf_vf_mux_scbd_156 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_156", this);
    pf_vf_mux_scbd_157 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_157", this);
    pf_vf_mux_scbd_158 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_158", this);
    pf_vf_mux_scbd_159 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_159", this);
    pf_vf_mux_scbd_160 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_160", this);
    pf_vf_mux_scbd_161 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_161", this);
    pf_vf_mux_scbd_162 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_162", this);
    pf_vf_mux_scbd_163 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_163", this);
    pf_vf_mux_scbd_164 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_164", this);
    pf_vf_mux_scbd_165 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_165", this);
    pf_vf_mux_scbd_166 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_166", this);
    pf_vf_mux_scbd_167 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_167", this);
    pf_vf_mux_scbd_168 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_168", this);
    pf_vf_mux_scbd_169 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_169", this);
    pf_vf_mux_scbd_170 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_170", this);
    pf_vf_mux_scbd_171 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_171", this);
    pf_vf_mux_scbd_172 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_172", this);
    pf_vf_mux_scbd_173 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_173", this);
    pf_vf_mux_scbd_174 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_174", this);
    pf_vf_mux_scbd_175 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_175", this);
    pf_vf_mux_scbd_176 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_176", this);
    pf_vf_mux_scbd_177 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_177", this);
    pf_vf_mux_scbd_178 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_178", this);
    pf_vf_mux_scbd_179 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_179", this);
    pf_vf_mux_scbd_180 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_180", this);
    pf_vf_mux_scbd_181 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_181", this);
    pf_vf_mux_scbd_182 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_182", this);
    pf_vf_mux_scbd_183 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_183", this);
    pf_vf_mux_scbd_184 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_184", this);
    pf_vf_mux_scbd_185 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_185", this);
    pf_vf_mux_scbd_186 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_186", this);
    pf_vf_mux_scbd_187 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_187", this);
    pf_vf_mux_scbd_188 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_188", this);
    pf_vf_mux_scbd_189 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_189", this);
    pf_vf_mux_scbd_190 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_190", this);
    pf_vf_mux_scbd_191 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_191", this);
    pf_vf_mux_scbd_192 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_192", this);
    pf_vf_mux_scbd_193 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_193", this);
    pf_vf_mux_scbd_194 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_194", this);
    pf_vf_mux_scbd_195 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_195", this);
    pf_vf_mux_scbd_196 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_196", this);
    pf_vf_mux_scbd_197 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_197", this);
    pf_vf_mux_scbd_198 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_198", this);
    pf_vf_mux_scbd_199 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_199", this);
    pf_vf_mux_scbd_200 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_200", this);
    pf_vf_mux_scbd_201 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_201", this);
    pf_vf_mux_scbd_202 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_202", this);
    pf_vf_mux_scbd_203 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_203", this);
    pf_vf_mux_scbd_204 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_204", this);
    pf_vf_mux_scbd_205 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_205", this);
    pf_vf_mux_scbd_206 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_206", this);
    pf_vf_mux_scbd_207 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_207", this);
    pf_vf_mux_scbd_208 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_208", this);
    pf_vf_mux_scbd_209 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_209", this);
    pf_vf_mux_scbd_210 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_210", this);
    pf_vf_mux_scbd_211 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_211", this);
    pf_vf_mux_scbd_212 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_212", this);
    pf_vf_mux_scbd_213 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_213", this);
    pf_vf_mux_scbd_214 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_214", this);
    pf_vf_mux_scbd_215 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_215", this);
    pf_vf_mux_scbd_216 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_216", this);
    pf_vf_mux_scbd_217 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_217", this);
    pf_vf_mux_scbd_218 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_218", this);
    pf_vf_mux_scbd_219 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_219", this);
    pf_vf_mux_scbd_220 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_220", this);
    pf_vf_mux_scbd_221 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_221", this);
    pf_vf_mux_scbd_222 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_222", this);
    pf_vf_mux_scbd_223 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_223", this);
    pf_vf_mux_scbd_224 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_224", this);
    pf_vf_mux_scbd_225 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_225", this);
    pf_vf_mux_scbd_226 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_226", this);
    pf_vf_mux_scbd_227 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_227", this);
    pf_vf_mux_scbd_228 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_228", this);
    pf_vf_mux_scbd_229 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_229", this);
    pf_vf_mux_scbd_230 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_230", this);
    pf_vf_mux_scbd_231 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_231", this);
    pf_vf_mux_scbd_232 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_232", this);
    pf_vf_mux_scbd_233 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_233", this);
    pf_vf_mux_scbd_234 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_234", this);
    pf_vf_mux_scbd_235 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_235", this);
    pf_vf_mux_scbd_236 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_236", this);
    pf_vf_mux_scbd_237 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_237", this);
    pf_vf_mux_scbd_238 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_238", this);
    pf_vf_mux_scbd_239 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_239", this);
    pf_vf_mux_scbd_240 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_240", this);
    pf_vf_mux_scbd_241 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_241", this);
    pf_vf_mux_scbd_242 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_242", this);
    pf_vf_mux_scbd_243 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_243", this);
    pf_vf_mux_scbd_244 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_244", this);
    pf_vf_mux_scbd_245 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_245", this);
    pf_vf_mux_scbd_246 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_246", this);
    pf_vf_mux_scbd_247 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_247", this);
    pf_vf_mux_scbd_248 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_248", this);
    pf_vf_mux_scbd_249 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_249", this);
    pf_vf_mux_scbd_250 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_250", this);
    pf_vf_mux_scbd_251 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_251", this);
    pf_vf_mux_scbd_252 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_252", this);
    pf_vf_mux_scbd_253 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_253", this);
    pf_vf_mux_scbd_254 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_254", this);
    pf_vf_mux_scbd_255 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_255", this);
    pf_vf_mux_scbd_256 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_256", this);
    pf_vf_mux_scbd_257 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_257", this);
    pf_vf_mux_scbd_258 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_258", this);
    pf_vf_mux_scbd_259 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_259", this);
    pf_vf_mux_scbd_260 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_260", this);
    pf_vf_mux_scbd_261 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_261", this);
    pf_vf_mux_scbd_262 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_262", this);
    pf_vf_mux_scbd_263 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_263", this);
    pf_vf_mux_scbd_264 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_264", this);
    pf_vf_mux_scbd_265 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_265", this);
    pf_vf_mux_scbd_266 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_266", this);
    pf_vf_mux_scbd_267 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_267", this);
    pf_vf_mux_scbd_268 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_268", this);
    pf_vf_mux_scbd_269 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_269", this);
    pf_vf_mux_scbd_270 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_270", this);
    pf_vf_mux_scbd_271 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_271", this);
    pf_vf_mux_scbd_272 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_272", this);
    pf_vf_mux_scbd_273 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_273", this);
    pf_vf_mux_scbd_274 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_274", this);
    pf_vf_mux_scbd_275 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_275", this);
    pf_vf_mux_scbd_276 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_276", this);
    pf_vf_mux_scbd_277 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_277", this);
    pf_vf_mux_scbd_278 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_278", this);
    pf_vf_mux_scbd_279 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_279", this);
    pf_vf_mux_scbd_280 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_280", this);
    pf_vf_mux_scbd_281 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_281", this);
    pf_vf_mux_scbd_282 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_282", this);
    pf_vf_mux_scbd_283 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_283", this);
    pf_vf_mux_scbd_284 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_284", this);
    pf_vf_mux_scbd_285 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_285", this);
    pf_vf_mux_scbd_286 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_286", this);
    pf_vf_mux_scbd_287 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_287", this);
    pf_vf_mux_scbd_288 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_288", this);
    pf_vf_mux_scbd_289 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_289", this);
    pf_vf_mux_scbd_290 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_290", this);
    pf_vf_mux_scbd_291 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_291", this);
    pf_vf_mux_scbd_292 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_292", this);
    pf_vf_mux_scbd_293 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_293", this);
    pf_vf_mux_scbd_294 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_294", this);
    pf_vf_mux_scbd_295 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_295", this);
    pf_vf_mux_scbd_296 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_296", this);
    pf_vf_mux_scbd_297 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_297", this);
    pf_vf_mux_scbd_298 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_298", this);
    pf_vf_mux_scbd_299 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_299", this);
    pf_vf_mux_scbd_300 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_300", this);
    pf_vf_mux_scbd_301 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_301", this);
    pf_vf_mux_scbd_302 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_302", this);
    pf_vf_mux_scbd_303 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_303", this);
    pf_vf_mux_scbd_304 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_304", this);
    pf_vf_mux_scbd_305 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_305", this);
    pf_vf_mux_scbd_306 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_306", this);
    pf_vf_mux_scbd_307 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_307", this);
    pf_vf_mux_scbd_308 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_308", this);
    pf_vf_mux_scbd_309 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_309", this);
    pf_vf_mux_scbd_310 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_310", this);
    pf_vf_mux_scbd_311 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_311", this);
    pf_vf_mux_scbd_312 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_312", this);
    pf_vf_mux_scbd_313 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_313", this);
    pf_vf_mux_scbd_314 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_314", this);
    pf_vf_mux_scbd_315 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_315", this);
    pf_vf_mux_scbd_316 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_316", this);
    pf_vf_mux_scbd_317 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_317", this);
    pf_vf_mux_scbd_318 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_318", this);
    pf_vf_mux_scbd_319 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_319", this);
    pf_vf_mux_scbd_320 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_320", this);
    pf_vf_mux_scbd_321 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_321", this);
    pf_vf_mux_scbd_322 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_322", this);
    pf_vf_mux_scbd_323 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_323", this);
    pf_vf_mux_scbd_324 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_324", this);
    pf_vf_mux_scbd_325 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_325", this);
    pf_vf_mux_scbd_326 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_326", this);
    pf_vf_mux_scbd_327 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_327", this);
    pf_vf_mux_scbd_328 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_328", this);
    pf_vf_mux_scbd_329 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_329", this);
    pf_vf_mux_scbd_330 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_330", this);
    pf_vf_mux_scbd_331 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_331", this);
    pf_vf_mux_scbd_332 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_332", this);
    pf_vf_mux_scbd_333 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_333", this);
    pf_vf_mux_scbd_334 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_334", this);
    pf_vf_mux_scbd_335 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_335", this);
    pf_vf_mux_scbd_336 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_336", this);
    pf_vf_mux_scbd_337 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_337", this);
    pf_vf_mux_scbd_338 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_338", this);
    pf_vf_mux_scbd_339 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_339", this);
    pf_vf_mux_scbd_340 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_340", this);
    pf_vf_mux_scbd_341 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_341", this);
    pf_vf_mux_scbd_342 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_342", this);
    pf_vf_mux_scbd_343 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_343", this);
    pf_vf_mux_scbd_344 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_344", this);
    pf_vf_mux_scbd_345 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_345", this);
    pf_vf_mux_scbd_346 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_346", this);
    pf_vf_mux_scbd_347 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_347", this);
    pf_vf_mux_scbd_348 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_348", this);
    pf_vf_mux_scbd_349 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_349", this);
    pf_vf_mux_scbd_350 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_350", this);
    pf_vf_mux_scbd_351 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_351", this);
    pf_vf_mux_scbd_352 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_352", this);
    pf_vf_mux_scbd_353 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_353", this);
    pf_vf_mux_scbd_354 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_354", this);
    pf_vf_mux_scbd_355 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_355", this);
    pf_vf_mux_scbd_356 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_356", this);
    pf_vf_mux_scbd_357 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_357", this);
    pf_vf_mux_scbd_358 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_358", this);
    pf_vf_mux_scbd_359 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_359", this);
    pf_vf_mux_scbd_360 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_360", this);
    pf_vf_mux_scbd_361 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_361", this);
    pf_vf_mux_scbd_362 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_362", this);
    pf_vf_mux_scbd_363 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_363", this);
    pf_vf_mux_scbd_364 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_364", this);
    pf_vf_mux_scbd_365 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_365", this);
    pf_vf_mux_scbd_366 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_366", this);
    pf_vf_mux_scbd_367 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_367", this);
    pf_vf_mux_scbd_368 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_368", this);
    pf_vf_mux_scbd_369 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_369", this);
    pf_vf_mux_scbd_370 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_370", this);
    pf_vf_mux_scbd_371 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_371", this);
    pf_vf_mux_scbd_372 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_372", this);
    pf_vf_mux_scbd_373 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_373", this);
    pf_vf_mux_scbd_374 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_374", this);
    pf_vf_mux_scbd_375 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_375", this);
    pf_vf_mux_scbd_376 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_376", this);
    pf_vf_mux_scbd_377 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_377", this);
    pf_vf_mux_scbd_378 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_378", this);
    pf_vf_mux_scbd_379 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_379", this);
    pf_vf_mux_scbd_380 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_380", this);
    pf_vf_mux_scbd_381 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_381", this);
    pf_vf_mux_scbd_382 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_382", this);
    pf_vf_mux_scbd_383 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_383", this);
    pf_vf_mux_scbd_384 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_384", this);
    pf_vf_mux_scbd_385 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_385", this);
    pf_vf_mux_scbd_386 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_386", this);
    pf_vf_mux_scbd_387 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_387", this);
    pf_vf_mux_scbd_388 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_388", this);
    pf_vf_mux_scbd_389 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_389", this);
    pf_vf_mux_scbd_390 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_390", this);
    pf_vf_mux_scbd_391 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_391", this);
    pf_vf_mux_scbd_392 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_392", this);
    pf_vf_mux_scbd_393 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_393", this);
    pf_vf_mux_scbd_394 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_394", this);
    pf_vf_mux_scbd_395 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_395", this);
    pf_vf_mux_scbd_396 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_396", this);
    pf_vf_mux_scbd_397 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_397", this);
    pf_vf_mux_scbd_398 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_398", this);
    pf_vf_mux_scbd_399 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_399", this);
    pf_vf_mux_scbd_400 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_400", this);
    pf_vf_mux_scbd_401 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_401", this);
    pf_vf_mux_scbd_402 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_402", this);
    pf_vf_mux_scbd_403 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_403", this);
    pf_vf_mux_scbd_404 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_404", this);
    pf_vf_mux_scbd_405 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_405", this);
    pf_vf_mux_scbd_406 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_406", this);
    pf_vf_mux_scbd_407 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_407", this);
    pf_vf_mux_scbd_408 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_408", this);
    pf_vf_mux_scbd_409 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_409", this);
    pf_vf_mux_scbd_410 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_410", this);
    pf_vf_mux_scbd_411 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_411", this);
    pf_vf_mux_scbd_412 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_412", this);
    pf_vf_mux_scbd_413 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_413", this);
    pf_vf_mux_scbd_414 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_414", this);
    pf_vf_mux_scbd_415 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_415", this);
    pf_vf_mux_scbd_416 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_416", this);
    pf_vf_mux_scbd_417 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_417", this);
    pf_vf_mux_scbd_418 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_418", this);
    pf_vf_mux_scbd_419 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_419", this);
    pf_vf_mux_scbd_420 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_420", this);
    pf_vf_mux_scbd_421 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_421", this);
    pf_vf_mux_scbd_422 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_422", this);
    pf_vf_mux_scbd_423 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_423", this);
    pf_vf_mux_scbd_424 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_424", this);
    pf_vf_mux_scbd_425 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_425", this);
    pf_vf_mux_scbd_426 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_426", this);
    pf_vf_mux_scbd_427 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_427", this);
    pf_vf_mux_scbd_428 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_428", this);
    pf_vf_mux_scbd_429 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_429", this);
    pf_vf_mux_scbd_430 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_430", this);
    pf_vf_mux_scbd_431 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_431", this);
    pf_vf_mux_scbd_432 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_432", this);
    pf_vf_mux_scbd_433 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_433", this);
    pf_vf_mux_scbd_434 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_434", this);
    pf_vf_mux_scbd_435 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_435", this);
    pf_vf_mux_scbd_436 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_436", this);
    pf_vf_mux_scbd_437 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_437", this);
    pf_vf_mux_scbd_438 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_438", this);
    pf_vf_mux_scbd_439 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_439", this);
    pf_vf_mux_scbd_440 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_440", this);
    pf_vf_mux_scbd_441 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_441", this);
    pf_vf_mux_scbd_442 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_442", this);
    pf_vf_mux_scbd_443 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_443", this);
    pf_vf_mux_scbd_444 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_444", this);
    pf_vf_mux_scbd_445 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_445", this);
    pf_vf_mux_scbd_446 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_446", this);
    pf_vf_mux_scbd_447 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_447", this);
    pf_vf_mux_scbd_448 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_448", this);
    pf_vf_mux_scbd_449 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_449", this);
    pf_vf_mux_scbd_450 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_450", this);
    pf_vf_mux_scbd_451 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_451", this);
    pf_vf_mux_scbd_452 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_452", this);
    pf_vf_mux_scbd_453 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_453", this);
    pf_vf_mux_scbd_454 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_454", this);
    pf_vf_mux_scbd_455 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_455", this);
    pf_vf_mux_scbd_456 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_456", this);
    pf_vf_mux_scbd_457 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_457", this);
    pf_vf_mux_scbd_458 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_458", this);
    pf_vf_mux_scbd_459 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_459", this);
    pf_vf_mux_scbd_460 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_460", this);
    pf_vf_mux_scbd_461 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_461", this);
    pf_vf_mux_scbd_462 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_462", this);
    pf_vf_mux_scbd_463 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_463", this);
    pf_vf_mux_scbd_464 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_464", this);
    pf_vf_mux_scbd_465 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_465", this);
    pf_vf_mux_scbd_466 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_466", this);
    pf_vf_mux_scbd_467 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_467", this);
    pf_vf_mux_scbd_468 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_468", this);
    pf_vf_mux_scbd_469 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_469", this);
    pf_vf_mux_scbd_470 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_470", this);
    pf_vf_mux_scbd_471 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_471", this);
    pf_vf_mux_scbd_472 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_472", this);
    pf_vf_mux_scbd_473 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_473", this);
    pf_vf_mux_scbd_474 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_474", this);
    pf_vf_mux_scbd_475 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_475", this);
    pf_vf_mux_scbd_476 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_476", this);
    pf_vf_mux_scbd_477 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_477", this);
    pf_vf_mux_scbd_478 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_478", this);
    pf_vf_mux_scbd_479 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_479", this);
    pf_vf_mux_scbd_480 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_480", this);
    pf_vf_mux_scbd_481 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_481", this);
    pf_vf_mux_scbd_482 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_482", this);
    pf_vf_mux_scbd_483 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_483", this);
    pf_vf_mux_scbd_484 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_484", this);
    pf_vf_mux_scbd_485 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_485", this);
    pf_vf_mux_scbd_486 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_486", this);
    pf_vf_mux_scbd_487 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_487", this);
    pf_vf_mux_scbd_488 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_488", this);
    pf_vf_mux_scbd_489 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_489", this);
    pf_vf_mux_scbd_490 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_490", this);
    pf_vf_mux_scbd_491 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_491", this);
    pf_vf_mux_scbd_492 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_492", this);
    pf_vf_mux_scbd_493 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_493", this);
    pf_vf_mux_scbd_494 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_494", this);
    pf_vf_mux_scbd_495 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_495", this);
    pf_vf_mux_scbd_496 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_496", this);
    pf_vf_mux_scbd_497 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_497", this);
    pf_vf_mux_scbd_498 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_498", this);
    pf_vf_mux_scbd_499 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_499", this);
    pf_vf_mux_scbd_500 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_500", this);
    pf_vf_mux_scbd_501 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_501", this);
    pf_vf_mux_scbd_502 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_502", this);
    pf_vf_mux_scbd_503 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_503", this);
    pf_vf_mux_scbd_504 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_504", this);
    pf_vf_mux_scbd_505 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_505", this);
    pf_vf_mux_scbd_506 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_506", this);
    pf_vf_mux_scbd_507 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_507", this);
    pf_vf_mux_scbd_508 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_508", this);
    pf_vf_mux_scbd_509 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_509", this);
    pf_vf_mux_scbd_510 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_510", this);
    pf_vf_mux_scbd_511 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_511", this);
    pf_vf_mux_scbd_512 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_512", this);
    pf_vf_mux_scbd_513 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_513", this);
    pf_vf_mux_scbd_514 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_514", this);
    pf_vf_mux_scbd_515 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_515", this);
    pf_vf_mux_scbd_516 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_516", this);
    pf_vf_mux_scbd_517 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_517", this);
    pf_vf_mux_scbd_518 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_518", this);
    pf_vf_mux_scbd_519 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_519", this);
    pf_vf_mux_scbd_520 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_520", this);
    pf_vf_mux_scbd_521 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_521", this);
    pf_vf_mux_scbd_522 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_522", this);
    pf_vf_mux_scbd_523 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_523", this);
    pf_vf_mux_scbd_524 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_524", this);
    pf_vf_mux_scbd_525 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_525", this);
    pf_vf_mux_scbd_526 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_526", this);
    pf_vf_mux_scbd_527 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_527", this);
    pf_vf_mux_scbd_528 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_528", this);
    pf_vf_mux_scbd_529 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_529", this);
    pf_vf_mux_scbd_530 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_530", this);
    pf_vf_mux_scbd_531 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_531", this);
    pf_vf_mux_scbd_532 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_532", this);
    pf_vf_mux_scbd_533 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_533", this);
    pf_vf_mux_scbd_534 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_534", this);
    pf_vf_mux_scbd_535 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_535", this);
    pf_vf_mux_scbd_536 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_536", this);
    pf_vf_mux_scbd_537 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_537", this);
    pf_vf_mux_scbd_538 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_538", this);
    pf_vf_mux_scbd_539 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_539", this);
    pf_vf_mux_scbd_540 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_540", this);
    pf_vf_mux_scbd_541 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_541", this);
    pf_vf_mux_scbd_542 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_542", this);
    pf_vf_mux_scbd_543 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_543", this);
    pf_vf_mux_scbd_544 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_544", this);
    pf_vf_mux_scbd_545 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_545", this);
    pf_vf_mux_scbd_546 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_546", this);
    pf_vf_mux_scbd_547 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_547", this);
    pf_vf_mux_scbd_548 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_548", this);
    pf_vf_mux_scbd_549 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_549", this);
    pf_vf_mux_scbd_550 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_550", this);
    pf_vf_mux_scbd_551 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_551", this);
    pf_vf_mux_scbd_552 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_552", this);
    pf_vf_mux_scbd_553 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_553", this);
    pf_vf_mux_scbd_554 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_554", this);
    pf_vf_mux_scbd_555 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_555", this);
    pf_vf_mux_scbd_556 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_556", this);
    pf_vf_mux_scbd_557 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_557", this);
    pf_vf_mux_scbd_558 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_558", this);
    pf_vf_mux_scbd_559 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_559", this);
    pf_vf_mux_scbd_560 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_560", this);
    pf_vf_mux_scbd_561 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_561", this);
    pf_vf_mux_scbd_562 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_562", this);
    pf_vf_mux_scbd_563 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_563", this);
    pf_vf_mux_scbd_564 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_564", this);
    pf_vf_mux_scbd_565 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_565", this);
    pf_vf_mux_scbd_566 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_566", this);
    pf_vf_mux_scbd_567 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_567", this);
    pf_vf_mux_scbd_568 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_568", this);
    pf_vf_mux_scbd_569 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_569", this);
    pf_vf_mux_scbd_570 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_570", this);
    pf_vf_mux_scbd_571 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_571", this);
    pf_vf_mux_scbd_572 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_572", this);
    pf_vf_mux_scbd_573 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_573", this);
    pf_vf_mux_scbd_574 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_574", this);
    pf_vf_mux_scbd_575 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_575", this);
    pf_vf_mux_scbd_576 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_576", this);
    pf_vf_mux_scbd_577 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_577", this);
    pf_vf_mux_scbd_578 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_578", this);
    pf_vf_mux_scbd_579 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_579", this);
    pf_vf_mux_scbd_580 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_580", this);
    pf_vf_mux_scbd_581 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_581", this);
    pf_vf_mux_scbd_582 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_582", this);
    pf_vf_mux_scbd_583 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_583", this);
    pf_vf_mux_scbd_584 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_584", this);
    pf_vf_mux_scbd_585 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_585", this);
    pf_vf_mux_scbd_586 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_586", this);
    pf_vf_mux_scbd_587 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_587", this);
    pf_vf_mux_scbd_588 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_588", this);
    pf_vf_mux_scbd_589 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_589", this);
    pf_vf_mux_scbd_590 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_590", this);
    pf_vf_mux_scbd_591 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_591", this);
    pf_vf_mux_scbd_592 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_592", this);
    pf_vf_mux_scbd_593 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_593", this);
    pf_vf_mux_scbd_594 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_594", this);
    pf_vf_mux_scbd_595 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_595", this);
    pf_vf_mux_scbd_596 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_596", this);
    pf_vf_mux_scbd_597 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_597", this);
    pf_vf_mux_scbd_598 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_598", this);
    pf_vf_mux_scbd_599 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_599", this);
    pf_vf_mux_scbd_600 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_600", this);
    pf_vf_mux_scbd_601 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_601", this);
    pf_vf_mux_scbd_602 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_602", this);
    pf_vf_mux_scbd_603 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_603", this);
    pf_vf_mux_scbd_604 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_604", this);
    pf_vf_mux_scbd_605 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_605", this);
    pf_vf_mux_scbd_606 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_606", this);
    pf_vf_mux_scbd_607 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_607", this);
    pf_vf_mux_scbd_608 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_608", this);
    pf_vf_mux_scbd_609 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_609", this);
    pf_vf_mux_scbd_610 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_610", this);
    pf_vf_mux_scbd_611 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_611", this);
    pf_vf_mux_scbd_612 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_612", this);
    pf_vf_mux_scbd_613 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_613", this);
    pf_vf_mux_scbd_614 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_614", this);
    pf_vf_mux_scbd_615 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_615", this);
    pf_vf_mux_scbd_616 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_616", this);
    pf_vf_mux_scbd_617 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_617", this);
    pf_vf_mux_scbd_618 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_618", this);
    pf_vf_mux_scbd_619 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_619", this);
    pf_vf_mux_scbd_620 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_620", this);
    pf_vf_mux_scbd_621 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_621", this);
    pf_vf_mux_scbd_622 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_622", this);
    pf_vf_mux_scbd_623 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_623", this);
    pf_vf_mux_scbd_624 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_624", this);
    pf_vf_mux_scbd_625 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_625", this);
    pf_vf_mux_scbd_626 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_626", this);
    pf_vf_mux_scbd_627 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_627", this);
    pf_vf_mux_scbd_628 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_628", this);
    pf_vf_mux_scbd_629 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_629", this);
    pf_vf_mux_scbd_630 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_630", this);
    pf_vf_mux_scbd_631 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_631", this);
    pf_vf_mux_scbd_632 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_632", this);
    pf_vf_mux_scbd_633 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_633", this);
    pf_vf_mux_scbd_634 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_634", this);
    pf_vf_mux_scbd_635 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_635", this);
    pf_vf_mux_scbd_636 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_636", this);
    pf_vf_mux_scbd_637 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_637", this);
    pf_vf_mux_scbd_638 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_638", this);
    pf_vf_mux_scbd_639 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_639", this);
    pf_vf_mux_scbd_640 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_640", this);
    pf_vf_mux_scbd_641 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_641", this);
    pf_vf_mux_scbd_642 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_642", this);
    pf_vf_mux_scbd_643 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_643", this);
    pf_vf_mux_scbd_644 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_644", this);
    pf_vf_mux_scbd_645 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_645", this);
    pf_vf_mux_scbd_646 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_646", this);
    pf_vf_mux_scbd_647 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_647", this);
    pf_vf_mux_scbd_648 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_648", this);
    pf_vf_mux_scbd_649 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_649", this);
    pf_vf_mux_scbd_650 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_650", this);
    pf_vf_mux_scbd_651 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_651", this);
    pf_vf_mux_scbd_652 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_652", this);
    pf_vf_mux_scbd_653 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_653", this);
    pf_vf_mux_scbd_654 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_654", this);
    pf_vf_mux_scbd_655 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_655", this);
    pf_vf_mux_scbd_656 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_656", this);
    pf_vf_mux_scbd_657 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_657", this);
    pf_vf_mux_scbd_658 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_658", this);
    pf_vf_mux_scbd_659 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_659", this);
    pf_vf_mux_scbd_660 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_660", this);
    pf_vf_mux_scbd_661 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_661", this);
    pf_vf_mux_scbd_662 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_662", this);
    pf_vf_mux_scbd_663 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_663", this);
    pf_vf_mux_scbd_664 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_664", this);
    pf_vf_mux_scbd_665 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_665", this);
    pf_vf_mux_scbd_666 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_666", this);
    pf_vf_mux_scbd_667 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_667", this);
    pf_vf_mux_scbd_668 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_668", this);
    pf_vf_mux_scbd_669 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_669", this);
    pf_vf_mux_scbd_670 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_670", this);
    pf_vf_mux_scbd_671 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_671", this);
    pf_vf_mux_scbd_672 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_672", this);
    pf_vf_mux_scbd_673 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_673", this);
    pf_vf_mux_scbd_674 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_674", this);
    pf_vf_mux_scbd_675 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_675", this);
    pf_vf_mux_scbd_676 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_676", this);
    pf_vf_mux_scbd_677 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_677", this);
    pf_vf_mux_scbd_678 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_678", this);
    pf_vf_mux_scbd_679 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_679", this);
    pf_vf_mux_scbd_680 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_680", this);
    pf_vf_mux_scbd_681 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_681", this);
    pf_vf_mux_scbd_682 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_682", this);
    pf_vf_mux_scbd_683 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_683", this);
    pf_vf_mux_scbd_684 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_684", this);
    pf_vf_mux_scbd_685 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_685", this);
    pf_vf_mux_scbd_686 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_686", this);
    pf_vf_mux_scbd_687 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_687", this);
    pf_vf_mux_scbd_688 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_688", this);
    pf_vf_mux_scbd_689 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_689", this);
    pf_vf_mux_scbd_690 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_690", this);
    pf_vf_mux_scbd_691 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_691", this);
    pf_vf_mux_scbd_692 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_692", this);
    pf_vf_mux_scbd_693 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_693", this);
    pf_vf_mux_scbd_694 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_694", this);
    pf_vf_mux_scbd_695 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_695", this);
    pf_vf_mux_scbd_696 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_696", this);
    pf_vf_mux_scbd_697 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_697", this);
    pf_vf_mux_scbd_698 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_698", this);
    pf_vf_mux_scbd_699 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_699", this);
    pf_vf_mux_scbd_700 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_700", this);
    pf_vf_mux_scbd_701 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_701", this);
    pf_vf_mux_scbd_702 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_702", this);
    pf_vf_mux_scbd_703 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_703", this);
    pf_vf_mux_scbd_704 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_704", this);
    pf_vf_mux_scbd_705 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_705", this);
    pf_vf_mux_scbd_706 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_706", this);
    pf_vf_mux_scbd_707 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_707", this);
    pf_vf_mux_scbd_708 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_708", this);
    pf_vf_mux_scbd_709 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_709", this);
    pf_vf_mux_scbd_710 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_710", this);
    pf_vf_mux_scbd_711 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_711", this);
    pf_vf_mux_scbd_712 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_712", this);
    pf_vf_mux_scbd_713 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_713", this);
    pf_vf_mux_scbd_714 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_714", this);
    pf_vf_mux_scbd_715 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_715", this);
    pf_vf_mux_scbd_716 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_716", this);
    pf_vf_mux_scbd_717 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_717", this);
    pf_vf_mux_scbd_718 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_718", this);
    pf_vf_mux_scbd_719 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_719", this);
    pf_vf_mux_scbd_720 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_720", this);
    pf_vf_mux_scbd_721 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_721", this);
    pf_vf_mux_scbd_722 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_722", this);
    pf_vf_mux_scbd_723 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_723", this);
    pf_vf_mux_scbd_724 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_724", this);
    pf_vf_mux_scbd_725 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_725", this);
    pf_vf_mux_scbd_726 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_726", this);
    pf_vf_mux_scbd_727 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_727", this);
    pf_vf_mux_scbd_728 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_728", this);
    pf_vf_mux_scbd_729 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_729", this);
    pf_vf_mux_scbd_730 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_730", this);
    pf_vf_mux_scbd_731 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_731", this);
    pf_vf_mux_scbd_732 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_732", this);
    pf_vf_mux_scbd_733 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_733", this);
    pf_vf_mux_scbd_734 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_734", this);
    pf_vf_mux_scbd_735 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_735", this);
    pf_vf_mux_scbd_736 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_736", this);
    pf_vf_mux_scbd_737 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_737", this);
    pf_vf_mux_scbd_738 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_738", this);
    pf_vf_mux_scbd_739 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_739", this);
    pf_vf_mux_scbd_740 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_740", this);
    pf_vf_mux_scbd_741 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_741", this);
    pf_vf_mux_scbd_742 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_742", this);
    pf_vf_mux_scbd_743 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_743", this);
    pf_vf_mux_scbd_744 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_744", this);
    pf_vf_mux_scbd_745 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_745", this);
    pf_vf_mux_scbd_746 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_746", this);
    pf_vf_mux_scbd_747 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_747", this);
    pf_vf_mux_scbd_748 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_748", this);
    pf_vf_mux_scbd_749 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_749", this);
    pf_vf_mux_scbd_750 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_750", this);
    pf_vf_mux_scbd_751 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_751", this);
    pf_vf_mux_scbd_752 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_752", this);
    pf_vf_mux_scbd_753 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_753", this);
    pf_vf_mux_scbd_754 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_754", this);
    pf_vf_mux_scbd_755 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_755", this);
    pf_vf_mux_scbd_756 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_756", this);
    pf_vf_mux_scbd_757 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_757", this);
    pf_vf_mux_scbd_758 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_758", this);
    pf_vf_mux_scbd_759 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_759", this);
    pf_vf_mux_scbd_760 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_760", this);
    pf_vf_mux_scbd_761 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_761", this);
    pf_vf_mux_scbd_762 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_762", this);
    pf_vf_mux_scbd_763 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_763", this);
    pf_vf_mux_scbd_764 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_764", this);
    pf_vf_mux_scbd_765 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_765", this);
    pf_vf_mux_scbd_766 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_766", this);
    pf_vf_mux_scbd_767 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_767", this);
    pf_vf_mux_scbd_768 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_768", this);
    pf_vf_mux_scbd_769 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_769", this);
    pf_vf_mux_scbd_770 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_770", this);
    pf_vf_mux_scbd_771 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_771", this);
    pf_vf_mux_scbd_772 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_772", this);
    pf_vf_mux_scbd_773 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_773", this);
    pf_vf_mux_scbd_774 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_774", this);
    pf_vf_mux_scbd_775 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_775", this);
    pf_vf_mux_scbd_776 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_776", this);
    pf_vf_mux_scbd_777 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_777", this);
    pf_vf_mux_scbd_778 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_778", this);
    pf_vf_mux_scbd_779 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_779", this);
    pf_vf_mux_scbd_780 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_780", this);
    pf_vf_mux_scbd_781 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_781", this);
    pf_vf_mux_scbd_782 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_782", this);
    pf_vf_mux_scbd_783 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_783", this);
    pf_vf_mux_scbd_784 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_784", this);
    pf_vf_mux_scbd_785 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_785", this);
    pf_vf_mux_scbd_786 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_786", this);
    pf_vf_mux_scbd_787 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_787", this);
    pf_vf_mux_scbd_788 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_788", this);
    pf_vf_mux_scbd_789 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_789", this);
    pf_vf_mux_scbd_790 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_790", this);
    pf_vf_mux_scbd_791 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_791", this);
    pf_vf_mux_scbd_792 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_792", this);
    pf_vf_mux_scbd_793 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_793", this);
    pf_vf_mux_scbd_794 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_794", this);
    pf_vf_mux_scbd_795 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_795", this);
    pf_vf_mux_scbd_796 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_796", this);
    pf_vf_mux_scbd_797 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_797", this);
    pf_vf_mux_scbd_798 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_798", this);
    pf_vf_mux_scbd_799 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_799", this);
    pf_vf_mux_scbd_800 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_800", this);
    pf_vf_mux_scbd_801 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_801", this);
    pf_vf_mux_scbd_802 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_802", this);
    pf_vf_mux_scbd_803 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_803", this);
    pf_vf_mux_scbd_804 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_804", this);
    pf_vf_mux_scbd_805 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_805", this);
    pf_vf_mux_scbd_806 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_806", this);
    pf_vf_mux_scbd_807 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_807", this);
    pf_vf_mux_scbd_808 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_808", this);
    pf_vf_mux_scbd_809 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_809", this);
    pf_vf_mux_scbd_810 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_810", this);
    pf_vf_mux_scbd_811 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_811", this);
    pf_vf_mux_scbd_812 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_812", this);
    pf_vf_mux_scbd_813 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_813", this);
    pf_vf_mux_scbd_814 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_814", this);
    pf_vf_mux_scbd_815 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_815", this);
    pf_vf_mux_scbd_816 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_816", this);
    pf_vf_mux_scbd_817 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_817", this);
    pf_vf_mux_scbd_818 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_818", this);
    pf_vf_mux_scbd_819 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_819", this);
    pf_vf_mux_scbd_820 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_820", this);
    pf_vf_mux_scbd_821 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_821", this);
    pf_vf_mux_scbd_822 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_822", this);
    pf_vf_mux_scbd_823 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_823", this);
    pf_vf_mux_scbd_824 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_824", this);
    pf_vf_mux_scbd_825 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_825", this);
    pf_vf_mux_scbd_826 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_826", this);
    pf_vf_mux_scbd_827 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_827", this);
    pf_vf_mux_scbd_828 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_828", this);
    pf_vf_mux_scbd_829 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_829", this);
    pf_vf_mux_scbd_830 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_830", this);
    pf_vf_mux_scbd_831 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_831", this);
    pf_vf_mux_scbd_832 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_832", this);
    pf_vf_mux_scbd_833 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_833", this);
    pf_vf_mux_scbd_834 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_834", this);
    pf_vf_mux_scbd_835 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_835", this);
    pf_vf_mux_scbd_836 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_836", this);
    pf_vf_mux_scbd_837 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_837", this);
    pf_vf_mux_scbd_838 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_838", this);
    pf_vf_mux_scbd_839 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_839", this);
    pf_vf_mux_scbd_840 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_840", this);
    pf_vf_mux_scbd_841 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_841", this);
    pf_vf_mux_scbd_842 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_842", this);
    pf_vf_mux_scbd_843 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_843", this);
    pf_vf_mux_scbd_844 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_844", this);
    pf_vf_mux_scbd_845 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_845", this);
    pf_vf_mux_scbd_846 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_846", this);
    pf_vf_mux_scbd_847 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_847", this);
    pf_vf_mux_scbd_848 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_848", this);
    pf_vf_mux_scbd_849 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_849", this);
    pf_vf_mux_scbd_850 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_850", this);
    pf_vf_mux_scbd_851 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_851", this);
    pf_vf_mux_scbd_852 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_852", this);
    pf_vf_mux_scbd_853 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_853", this);
    pf_vf_mux_scbd_854 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_854", this);
    pf_vf_mux_scbd_855 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_855", this);
    pf_vf_mux_scbd_856 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_856", this);
    pf_vf_mux_scbd_857 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_857", this);
    pf_vf_mux_scbd_858 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_858", this);
    pf_vf_mux_scbd_859 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_859", this);
    pf_vf_mux_scbd_860 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_860", this);
    pf_vf_mux_scbd_861 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_861", this);
    pf_vf_mux_scbd_862 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_862", this);
    pf_vf_mux_scbd_863 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_863", this);
    pf_vf_mux_scbd_864 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_864", this);
    pf_vf_mux_scbd_865 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_865", this);
    pf_vf_mux_scbd_866 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_866", this);
    pf_vf_mux_scbd_867 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_867", this);
    pf_vf_mux_scbd_868 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_868", this);
    pf_vf_mux_scbd_869 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_869", this);
    pf_vf_mux_scbd_870 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_870", this);
    pf_vf_mux_scbd_871 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_871", this);
    pf_vf_mux_scbd_872 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_872", this);
    pf_vf_mux_scbd_873 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_873", this);
    pf_vf_mux_scbd_874 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_874", this);
    pf_vf_mux_scbd_875 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_875", this);
    pf_vf_mux_scbd_876 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_876", this);
    pf_vf_mux_scbd_877 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_877", this);
    pf_vf_mux_scbd_878 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_878", this);
    pf_vf_mux_scbd_879 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_879", this);
    pf_vf_mux_scbd_880 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_880", this);
    pf_vf_mux_scbd_881 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_881", this);
    pf_vf_mux_scbd_882 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_882", this);
    pf_vf_mux_scbd_883 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_883", this);
    pf_vf_mux_scbd_884 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_884", this);
    pf_vf_mux_scbd_885 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_885", this);
    pf_vf_mux_scbd_886 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_886", this);
    pf_vf_mux_scbd_887 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_887", this);
    pf_vf_mux_scbd_888 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_888", this);
    pf_vf_mux_scbd_889 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_889", this);
    pf_vf_mux_scbd_890 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_890", this);
    pf_vf_mux_scbd_891 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_891", this);
    pf_vf_mux_scbd_892 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_892", this);
    pf_vf_mux_scbd_893 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_893", this);
    pf_vf_mux_scbd_894 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_894", this);
    pf_vf_mux_scbd_895 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_895", this);
    pf_vf_mux_scbd_896 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_896", this);
    pf_vf_mux_scbd_897 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_897", this);
    pf_vf_mux_scbd_898 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_898", this);
    pf_vf_mux_scbd_899 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_899", this);
    pf_vf_mux_scbd_900 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_900", this);
    pf_vf_mux_scbd_901 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_901", this);
    pf_vf_mux_scbd_902 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_902", this);
    pf_vf_mux_scbd_903 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_903", this);
    pf_vf_mux_scbd_904 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_904", this);
    pf_vf_mux_scbd_905 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_905", this);
    pf_vf_mux_scbd_906 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_906", this);
    pf_vf_mux_scbd_907 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_907", this);
    pf_vf_mux_scbd_908 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_908", this);
    pf_vf_mux_scbd_909 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_909", this);
    pf_vf_mux_scbd_910 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_910", this);
    pf_vf_mux_scbd_911 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_911", this);
    pf_vf_mux_scbd_912 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_912", this);
    pf_vf_mux_scbd_913 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_913", this);
    pf_vf_mux_scbd_914 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_914", this);
    pf_vf_mux_scbd_915 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_915", this);
    pf_vf_mux_scbd_916 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_916", this);
    pf_vf_mux_scbd_917 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_917", this);
    pf_vf_mux_scbd_918 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_918", this);
    pf_vf_mux_scbd_919 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_919", this);
    pf_vf_mux_scbd_920 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_920", this);
    pf_vf_mux_scbd_921 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_921", this);
    pf_vf_mux_scbd_922 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_922", this);
    pf_vf_mux_scbd_923 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_923", this);
    pf_vf_mux_scbd_924 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_924", this);
    pf_vf_mux_scbd_925 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_925", this);
    pf_vf_mux_scbd_926 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_926", this);
    pf_vf_mux_scbd_927 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_927", this);
    pf_vf_mux_scbd_928 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_928", this);
    pf_vf_mux_scbd_929 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_929", this);
    pf_vf_mux_scbd_930 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_930", this);
    pf_vf_mux_scbd_931 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_931", this);
    pf_vf_mux_scbd_932 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_932", this);
    pf_vf_mux_scbd_933 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_933", this);
    pf_vf_mux_scbd_934 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_934", this);
    pf_vf_mux_scbd_935 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_935", this);
    pf_vf_mux_scbd_936 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_936", this);
    pf_vf_mux_scbd_937 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_937", this);
    pf_vf_mux_scbd_938 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_938", this);
    pf_vf_mux_scbd_939 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_939", this);
    pf_vf_mux_scbd_940 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_940", this);
    pf_vf_mux_scbd_941 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_941", this);
    pf_vf_mux_scbd_942 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_942", this);
    pf_vf_mux_scbd_943 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_943", this);
    pf_vf_mux_scbd_944 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_944", this);
    pf_vf_mux_scbd_945 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_945", this);
    pf_vf_mux_scbd_946 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_946", this);
    pf_vf_mux_scbd_947 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_947", this);
    pf_vf_mux_scbd_948 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_948", this);
    pf_vf_mux_scbd_949 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_949", this);
    pf_vf_mux_scbd_950 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_950", this);
    pf_vf_mux_scbd_951 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_951", this);
    pf_vf_mux_scbd_952 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_952", this);
    pf_vf_mux_scbd_953 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_953", this);
    pf_vf_mux_scbd_954 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_954", this);
    pf_vf_mux_scbd_955 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_955", this);
    pf_vf_mux_scbd_956 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_956", this);
    pf_vf_mux_scbd_957 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_957", this);
    pf_vf_mux_scbd_958 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_958", this);
    pf_vf_mux_scbd_959 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_959", this);
    pf_vf_mux_scbd_960 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_960", this);
    pf_vf_mux_scbd_961 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_961", this);
    pf_vf_mux_scbd_962 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_962", this);
    pf_vf_mux_scbd_963 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_963", this);
    pf_vf_mux_scbd_964 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_964", this);
    pf_vf_mux_scbd_965 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_965", this);
    pf_vf_mux_scbd_966 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_966", this);
    pf_vf_mux_scbd_967 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_967", this);
    pf_vf_mux_scbd_968 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_968", this);
    pf_vf_mux_scbd_969 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_969", this);
    pf_vf_mux_scbd_970 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_970", this);
    pf_vf_mux_scbd_971 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_971", this);
    pf_vf_mux_scbd_972 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_972", this);
    pf_vf_mux_scbd_973 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_973", this);
    pf_vf_mux_scbd_974 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_974", this);
    pf_vf_mux_scbd_975 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_975", this);
    pf_vf_mux_scbd_976 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_976", this);
    pf_vf_mux_scbd_977 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_977", this);
    pf_vf_mux_scbd_978 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_978", this);
    pf_vf_mux_scbd_979 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_979", this);
    pf_vf_mux_scbd_980 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_980", this);
    pf_vf_mux_scbd_981 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_981", this);
    pf_vf_mux_scbd_982 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_982", this);
    pf_vf_mux_scbd_983 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_983", this);
    pf_vf_mux_scbd_984 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_984", this);
    pf_vf_mux_scbd_985 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_985", this);
    pf_vf_mux_scbd_986 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_986", this);
    pf_vf_mux_scbd_987 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_987", this);
    pf_vf_mux_scbd_988 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_988", this);
    pf_vf_mux_scbd_989 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_989", this);
    pf_vf_mux_scbd_990 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_990", this);
    pf_vf_mux_scbd_991 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_991", this);
    pf_vf_mux_scbd_992 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_992", this);
    pf_vf_mux_scbd_993 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_993", this);
    pf_vf_mux_scbd_994 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_994", this);
    pf_vf_mux_scbd_995 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_995", this);
    pf_vf_mux_scbd_996 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_996", this);
    pf_vf_mux_scbd_997 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_997", this);
    pf_vf_mux_scbd_998 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_998", this);
    pf_vf_mux_scbd_999 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_999", this);
    pf_vf_mux_scbd_1000 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1000", this);
    pf_vf_mux_scbd_1001 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1001", this);
    pf_vf_mux_scbd_1002 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1002", this);
    pf_vf_mux_scbd_1003 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1003", this);
    pf_vf_mux_scbd_1004 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1004", this);
    pf_vf_mux_scbd_1005 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1005", this);
    pf_vf_mux_scbd_1006 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1006", this);
    pf_vf_mux_scbd_1007 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1007", this);
    pf_vf_mux_scbd_1008 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1008", this);
    pf_vf_mux_scbd_1009 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1009", this);
    pf_vf_mux_scbd_1010 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1010", this);
    pf_vf_mux_scbd_1011 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1011", this);
    pf_vf_mux_scbd_1012 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1012", this);
    pf_vf_mux_scbd_1013 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1013", this);
    pf_vf_mux_scbd_1014 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1014", this);
    pf_vf_mux_scbd_1015 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1015", this);
    pf_vf_mux_scbd_1016 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1016", this);
    pf_vf_mux_scbd_1017 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1017", this);
    pf_vf_mux_scbd_1018 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1018", this);
    pf_vf_mux_scbd_1019 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1019", this);
    pf_vf_mux_scbd_1020 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1020", this);
    pf_vf_mux_scbd_1021 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1021", this);
    pf_vf_mux_scbd_1022 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1022", this);
    pf_vf_mux_scbd_1023 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1023", this);
    pf_vf_mux_scbd_1024 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1024", this);
    pf_vf_mux_scbd_1025 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1025", this);
    pf_vf_mux_scbd_1026 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1026", this);
    pf_vf_mux_scbd_1027 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1027", this);
    pf_vf_mux_scbd_1028 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1028", this);
    pf_vf_mux_scbd_1029 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1029", this);
    pf_vf_mux_scbd_1030 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1030", this);
    pf_vf_mux_scbd_1031 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1031", this);
    pf_vf_mux_scbd_1032 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1032", this);
    pf_vf_mux_scbd_1033 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1033", this);
    pf_vf_mux_scbd_1034 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1034", this);
    pf_vf_mux_scbd_1035 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1035", this);
    pf_vf_mux_scbd_1036 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1036", this);
    pf_vf_mux_scbd_1037 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1037", this);
    pf_vf_mux_scbd_1038 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1038", this);
    pf_vf_mux_scbd_1039 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1039", this);
    pf_vf_mux_scbd_1040 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1040", this);
    pf_vf_mux_scbd_1041 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1041", this);
    pf_vf_mux_scbd_1042 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1042", this);
    pf_vf_mux_scbd_1043 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1043", this);
    pf_vf_mux_scbd_1044 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1044", this);
    pf_vf_mux_scbd_1045 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1045", this);
    pf_vf_mux_scbd_1046 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1046", this);
    pf_vf_mux_scbd_1047 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1047", this);
    pf_vf_mux_scbd_1048 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1048", this);
    pf_vf_mux_scbd_1049 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1049", this);
    pf_vf_mux_scbd_1050 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1050", this);
    pf_vf_mux_scbd_1051 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1051", this);
    pf_vf_mux_scbd_1052 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1052", this);
    pf_vf_mux_scbd_1053 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1053", this);
    pf_vf_mux_scbd_1054 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1054", this);
    pf_vf_mux_scbd_1055 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1055", this);
    pf_vf_mux_scbd_1056 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1056", this);
    pf_vf_mux_scbd_1057 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1057", this);
    pf_vf_mux_scbd_1058 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1058", this);
    pf_vf_mux_scbd_1059 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1059", this);
    pf_vf_mux_scbd_1060 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1060", this);
    pf_vf_mux_scbd_1061 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1061", this);
    pf_vf_mux_scbd_1062 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1062", this);
    pf_vf_mux_scbd_1063 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1063", this);
    pf_vf_mux_scbd_1064 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1064", this);
    pf_vf_mux_scbd_1065 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1065", this);
    pf_vf_mux_scbd_1066 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1066", this);
    pf_vf_mux_scbd_1067 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1067", this);
    pf_vf_mux_scbd_1068 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1068", this);
    pf_vf_mux_scbd_1069 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1069", this);
    pf_vf_mux_scbd_1070 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1070", this);
    pf_vf_mux_scbd_1071 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1071", this);
    pf_vf_mux_scbd_1072 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1072", this);
    pf_vf_mux_scbd_1073 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1073", this);
    pf_vf_mux_scbd_1074 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1074", this);
    pf_vf_mux_scbd_1075 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1075", this);
    pf_vf_mux_scbd_1076 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1076", this);
    pf_vf_mux_scbd_1077 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1077", this);
    pf_vf_mux_scbd_1078 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1078", this);
    pf_vf_mux_scbd_1079 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1079", this);
    pf_vf_mux_scbd_1080 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1080", this);
    pf_vf_mux_scbd_1081 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1081", this);
    pf_vf_mux_scbd_1082 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1082", this);
    pf_vf_mux_scbd_1083 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1083", this);
    pf_vf_mux_scbd_1084 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1084", this);
    pf_vf_mux_scbd_1085 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1085", this);
    pf_vf_mux_scbd_1086 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1086", this);
    pf_vf_mux_scbd_1087 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1087", this);
    pf_vf_mux_scbd_1088 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1088", this);
    pf_vf_mux_scbd_1089 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1089", this);
    pf_vf_mux_scbd_1090 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1090", this);
    pf_vf_mux_scbd_1091 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1091", this);
    pf_vf_mux_scbd_1092 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1092", this);
    pf_vf_mux_scbd_1093 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1093", this);
    pf_vf_mux_scbd_1094 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1094", this);
    pf_vf_mux_scbd_1095 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1095", this);
    pf_vf_mux_scbd_1096 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1096", this);
    pf_vf_mux_scbd_1097 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1097", this);
    pf_vf_mux_scbd_1098 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1098", this);
    pf_vf_mux_scbd_1099 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1099", this);
    pf_vf_mux_scbd_1100 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1100", this);
    pf_vf_mux_scbd_1101 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1101", this);
    pf_vf_mux_scbd_1102 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1102", this);
    pf_vf_mux_scbd_1103 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1103", this);
    pf_vf_mux_scbd_1104 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1104", this);
    pf_vf_mux_scbd_1105 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1105", this);
    pf_vf_mux_scbd_1106 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1106", this);
    pf_vf_mux_scbd_1107 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1107", this);
    pf_vf_mux_scbd_1108 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1108", this);
    pf_vf_mux_scbd_1109 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1109", this);
    pf_vf_mux_scbd_1110 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1110", this);
    pf_vf_mux_scbd_1111 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1111", this);
    pf_vf_mux_scbd_1112 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1112", this);
    pf_vf_mux_scbd_1113 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1113", this);
    pf_vf_mux_scbd_1114 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1114", this);
    pf_vf_mux_scbd_1115 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1115", this);
    pf_vf_mux_scbd_1116 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1116", this);
    pf_vf_mux_scbd_1117 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1117", this);
    pf_vf_mux_scbd_1118 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1118", this);
    pf_vf_mux_scbd_1119 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1119", this);
    pf_vf_mux_scbd_1120 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1120", this);
    pf_vf_mux_scbd_1121 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1121", this);
    pf_vf_mux_scbd_1122 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1122", this);
    pf_vf_mux_scbd_1123 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1123", this);
    pf_vf_mux_scbd_1124 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1124", this);
    pf_vf_mux_scbd_1125 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1125", this);
    pf_vf_mux_scbd_1126 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1126", this);
    pf_vf_mux_scbd_1127 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1127", this);
    pf_vf_mux_scbd_1128 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1128", this);
    pf_vf_mux_scbd_1129 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1129", this);
    pf_vf_mux_scbd_1130 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1130", this);
    pf_vf_mux_scbd_1131 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1131", this);
    pf_vf_mux_scbd_1132 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1132", this);
    pf_vf_mux_scbd_1133 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1133", this);
    pf_vf_mux_scbd_1134 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1134", this);
    pf_vf_mux_scbd_1135 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1135", this);
    pf_vf_mux_scbd_1136 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1136", this);
    pf_vf_mux_scbd_1137 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1137", this);
    pf_vf_mux_scbd_1138 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1138", this);
    pf_vf_mux_scbd_1139 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1139", this);
    pf_vf_mux_scbd_1140 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1140", this);
    pf_vf_mux_scbd_1141 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1141", this);
    pf_vf_mux_scbd_1142 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1142", this);
    pf_vf_mux_scbd_1143 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1143", this);
    pf_vf_mux_scbd_1144 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1144", this);
    pf_vf_mux_scbd_1145 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1145", this);
    pf_vf_mux_scbd_1146 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1146", this);
    pf_vf_mux_scbd_1147 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1147", this);
    pf_vf_mux_scbd_1148 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1148", this);
    pf_vf_mux_scbd_1149 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1149", this);
    pf_vf_mux_scbd_1150 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1150", this);
    pf_vf_mux_scbd_1151 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1151", this);
    pf_vf_mux_scbd_1152 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1152", this);
    pf_vf_mux_scbd_1153 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1153", this);
    pf_vf_mux_scbd_1154 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1154", this);
    pf_vf_mux_scbd_1155 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1155", this);
    pf_vf_mux_scbd_1156 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1156", this);
    pf_vf_mux_scbd_1157 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1157", this);
    pf_vf_mux_scbd_1158 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1158", this);
    pf_vf_mux_scbd_1159 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1159", this);
    pf_vf_mux_scbd_1160 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1160", this);
    pf_vf_mux_scbd_1161 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1161", this);
    pf_vf_mux_scbd_1162 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1162", this);
    pf_vf_mux_scbd_1163 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1163", this);
    pf_vf_mux_scbd_1164 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1164", this);
    pf_vf_mux_scbd_1165 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1165", this);
    pf_vf_mux_scbd_1166 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1166", this);
    pf_vf_mux_scbd_1167 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1167", this);
    pf_vf_mux_scbd_1168 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1168", this);
    pf_vf_mux_scbd_1169 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1169", this);
    pf_vf_mux_scbd_1170 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1170", this);
    pf_vf_mux_scbd_1171 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1171", this);
    pf_vf_mux_scbd_1172 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1172", this);
    pf_vf_mux_scbd_1173 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1173", this);
    pf_vf_mux_scbd_1174 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1174", this);
    pf_vf_mux_scbd_1175 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1175", this);
    pf_vf_mux_scbd_1176 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1176", this);
    pf_vf_mux_scbd_1177 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1177", this);
    pf_vf_mux_scbd_1178 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1178", this);
    pf_vf_mux_scbd_1179 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1179", this);
    pf_vf_mux_scbd_1180 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1180", this);
    pf_vf_mux_scbd_1181 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1181", this);
    pf_vf_mux_scbd_1182 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1182", this);
    pf_vf_mux_scbd_1183 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1183", this);
    pf_vf_mux_scbd_1184 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1184", this);
    pf_vf_mux_scbd_1185 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1185", this);
    pf_vf_mux_scbd_1186 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1186", this);
    pf_vf_mux_scbd_1187 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1187", this);
    pf_vf_mux_scbd_1188 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1188", this);
    pf_vf_mux_scbd_1189 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1189", this);
    pf_vf_mux_scbd_1190 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1190", this);
    pf_vf_mux_scbd_1191 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1191", this);
    pf_vf_mux_scbd_1192 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1192", this);
    pf_vf_mux_scbd_1193 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1193", this);
    pf_vf_mux_scbd_1194 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1194", this);
    pf_vf_mux_scbd_1195 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1195", this);
    pf_vf_mux_scbd_1196 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1196", this);
    pf_vf_mux_scbd_1197 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1197", this);
    pf_vf_mux_scbd_1198 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1198", this);
    pf_vf_mux_scbd_1199 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1199", this);
    pf_vf_mux_scbd_1200 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1200", this);
    pf_vf_mux_scbd_1201 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1201", this);
    pf_vf_mux_scbd_1202 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1202", this);
    pf_vf_mux_scbd_1203 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1203", this);
    pf_vf_mux_scbd_1204 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1204", this);
    pf_vf_mux_scbd_1205 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1205", this);
    pf_vf_mux_scbd_1206 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1206", this);
    pf_vf_mux_scbd_1207 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1207", this);
    pf_vf_mux_scbd_1208 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1208", this);
    pf_vf_mux_scbd_1209 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1209", this);
    pf_vf_mux_scbd_1210 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1210", this);
    pf_vf_mux_scbd_1211 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1211", this);
    pf_vf_mux_scbd_1212 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1212", this);
    pf_vf_mux_scbd_1213 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1213", this);
    pf_vf_mux_scbd_1214 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1214", this);
    pf_vf_mux_scbd_1215 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1215", this);
    pf_vf_mux_scbd_1216 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1216", this);
    pf_vf_mux_scbd_1217 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1217", this);
    pf_vf_mux_scbd_1218 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1218", this);
    pf_vf_mux_scbd_1219 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1219", this);
    pf_vf_mux_scbd_1220 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1220", this);
    pf_vf_mux_scbd_1221 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1221", this);
    pf_vf_mux_scbd_1222 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1222", this);
    pf_vf_mux_scbd_1223 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1223", this);
    pf_vf_mux_scbd_1224 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1224", this);
    pf_vf_mux_scbd_1225 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1225", this);
    pf_vf_mux_scbd_1226 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1226", this);
    pf_vf_mux_scbd_1227 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1227", this);
    pf_vf_mux_scbd_1228 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1228", this);
    pf_vf_mux_scbd_1229 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1229", this);
    pf_vf_mux_scbd_1230 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1230", this);
    pf_vf_mux_scbd_1231 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1231", this);
    pf_vf_mux_scbd_1232 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1232", this);
    pf_vf_mux_scbd_1233 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1233", this);
    pf_vf_mux_scbd_1234 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1234", this);
    pf_vf_mux_scbd_1235 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1235", this);
    pf_vf_mux_scbd_1236 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1236", this);
    pf_vf_mux_scbd_1237 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1237", this);
    pf_vf_mux_scbd_1238 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1238", this);
    pf_vf_mux_scbd_1239 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1239", this);
    pf_vf_mux_scbd_1240 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1240", this);
    pf_vf_mux_scbd_1241 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1241", this);
    pf_vf_mux_scbd_1242 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1242", this);
    pf_vf_mux_scbd_1243 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1243", this);
    pf_vf_mux_scbd_1244 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1244", this);
    pf_vf_mux_scbd_1245 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1245", this);
    pf_vf_mux_scbd_1246 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1246", this);
    pf_vf_mux_scbd_1247 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1247", this);
    pf_vf_mux_scbd_1248 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1248", this);
    pf_vf_mux_scbd_1249 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1249", this);
    pf_vf_mux_scbd_1250 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1250", this);
    pf_vf_mux_scbd_1251 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1251", this);
    pf_vf_mux_scbd_1252 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1252", this);
    pf_vf_mux_scbd_1253 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1253", this);
    pf_vf_mux_scbd_1254 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1254", this);
    pf_vf_mux_scbd_1255 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1255", this);
    pf_vf_mux_scbd_1256 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1256", this);
    pf_vf_mux_scbd_1257 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1257", this);
    pf_vf_mux_scbd_1258 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1258", this);
    pf_vf_mux_scbd_1259 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1259", this);
    pf_vf_mux_scbd_1260 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1260", this);
    pf_vf_mux_scbd_1261 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1261", this);
    pf_vf_mux_scbd_1262 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1262", this);
    pf_vf_mux_scbd_1263 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1263", this);
    pf_vf_mux_scbd_1264 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1264", this);
    pf_vf_mux_scbd_1265 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1265", this);
    pf_vf_mux_scbd_1266 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1266", this);
    pf_vf_mux_scbd_1267 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1267", this);
    pf_vf_mux_scbd_1268 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1268", this);
    pf_vf_mux_scbd_1269 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1269", this);
    pf_vf_mux_scbd_1270 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1270", this);
    pf_vf_mux_scbd_1271 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1271", this);
    pf_vf_mux_scbd_1272 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1272", this);
    pf_vf_mux_scbd_1273 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1273", this);
    pf_vf_mux_scbd_1274 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1274", this);
    pf_vf_mux_scbd_1275 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1275", this);
    pf_vf_mux_scbd_1276 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1276", this);
    pf_vf_mux_scbd_1277 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1277", this);
    pf_vf_mux_scbd_1278 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1278", this);
    pf_vf_mux_scbd_1279 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1279", this);
    pf_vf_mux_scbd_1280 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1280", this);
    pf_vf_mux_scbd_1281 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1281", this);
    pf_vf_mux_scbd_1282 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1282", this);
    pf_vf_mux_scbd_1283 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1283", this);
    pf_vf_mux_scbd_1284 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1284", this);
    pf_vf_mux_scbd_1285 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1285", this);
    pf_vf_mux_scbd_1286 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1286", this);
    pf_vf_mux_scbd_1287 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1287", this);
    pf_vf_mux_scbd_1288 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1288", this);
    pf_vf_mux_scbd_1289 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1289", this);
    pf_vf_mux_scbd_1290 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1290", this);
    pf_vf_mux_scbd_1291 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1291", this);
    pf_vf_mux_scbd_1292 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1292", this);
    pf_vf_mux_scbd_1293 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1293", this);
    pf_vf_mux_scbd_1294 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1294", this);
    pf_vf_mux_scbd_1295 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1295", this);
    pf_vf_mux_scbd_1296 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1296", this);
    pf_vf_mux_scbd_1297 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1297", this);
    pf_vf_mux_scbd_1298 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1298", this);
    pf_vf_mux_scbd_1299 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1299", this);
    pf_vf_mux_scbd_1300 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1300", this);
    pf_vf_mux_scbd_1301 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1301", this);
    pf_vf_mux_scbd_1302 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1302", this);
    pf_vf_mux_scbd_1303 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1303", this);
    pf_vf_mux_scbd_1304 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1304", this);
    pf_vf_mux_scbd_1305 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1305", this);
    pf_vf_mux_scbd_1306 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1306", this);
    pf_vf_mux_scbd_1307 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1307", this);
    pf_vf_mux_scbd_1308 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1308", this);
    pf_vf_mux_scbd_1309 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1309", this);
    pf_vf_mux_scbd_1310 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1310", this);
    pf_vf_mux_scbd_1311 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1311", this);
    pf_vf_mux_scbd_1312 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1312", this);
    pf_vf_mux_scbd_1313 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1313", this);
    pf_vf_mux_scbd_1314 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1314", this);
    pf_vf_mux_scbd_1315 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1315", this);
    pf_vf_mux_scbd_1316 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1316", this);
    pf_vf_mux_scbd_1317 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1317", this);
    pf_vf_mux_scbd_1318 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1318", this);
    pf_vf_mux_scbd_1319 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1319", this);
    pf_vf_mux_scbd_1320 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1320", this);
    pf_vf_mux_scbd_1321 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1321", this);
    pf_vf_mux_scbd_1322 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1322", this);
    pf_vf_mux_scbd_1323 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1323", this);
    pf_vf_mux_scbd_1324 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1324", this);
    pf_vf_mux_scbd_1325 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1325", this);
    pf_vf_mux_scbd_1326 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1326", this);
    pf_vf_mux_scbd_1327 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1327", this);
    pf_vf_mux_scbd_1328 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1328", this);
    pf_vf_mux_scbd_1329 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1329", this);
    pf_vf_mux_scbd_1330 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1330", this);
    pf_vf_mux_scbd_1331 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1331", this);
    pf_vf_mux_scbd_1332 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1332", this);
    pf_vf_mux_scbd_1333 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1333", this);
    pf_vf_mux_scbd_1334 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1334", this);
    pf_vf_mux_scbd_1335 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1335", this);
    pf_vf_mux_scbd_1336 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1336", this);
    pf_vf_mux_scbd_1337 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1337", this);
    pf_vf_mux_scbd_1338 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1338", this);
    pf_vf_mux_scbd_1339 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1339", this);
    pf_vf_mux_scbd_1340 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1340", this);
    pf_vf_mux_scbd_1341 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1341", this);
    pf_vf_mux_scbd_1342 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1342", this);
    pf_vf_mux_scbd_1343 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1343", this);
    pf_vf_mux_scbd_1344 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1344", this);
    pf_vf_mux_scbd_1345 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1345", this);
    pf_vf_mux_scbd_1346 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1346", this);
    pf_vf_mux_scbd_1347 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1347", this);
    pf_vf_mux_scbd_1348 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1348", this);
    pf_vf_mux_scbd_1349 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1349", this);
    pf_vf_mux_scbd_1350 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1350", this);
    pf_vf_mux_scbd_1351 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1351", this);
    pf_vf_mux_scbd_1352 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1352", this);
    pf_vf_mux_scbd_1353 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1353", this);
    pf_vf_mux_scbd_1354 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1354", this);
    pf_vf_mux_scbd_1355 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1355", this);
    pf_vf_mux_scbd_1356 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1356", this);
    pf_vf_mux_scbd_1357 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1357", this);
    pf_vf_mux_scbd_1358 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1358", this);
    pf_vf_mux_scbd_1359 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1359", this);
    pf_vf_mux_scbd_1360 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1360", this);
    pf_vf_mux_scbd_1361 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1361", this);
    pf_vf_mux_scbd_1362 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1362", this);
    pf_vf_mux_scbd_1363 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1363", this);
    pf_vf_mux_scbd_1364 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1364", this);
    pf_vf_mux_scbd_1365 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1365", this);
    pf_vf_mux_scbd_1366 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1366", this);
    pf_vf_mux_scbd_1367 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1367", this);
    pf_vf_mux_scbd_1368 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1368", this);
    pf_vf_mux_scbd_1369 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1369", this);
    pf_vf_mux_scbd_1370 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1370", this);
    pf_vf_mux_scbd_1371 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1371", this);
    pf_vf_mux_scbd_1372 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1372", this);
    pf_vf_mux_scbd_1373 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1373", this);
    pf_vf_mux_scbd_1374 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1374", this);
    pf_vf_mux_scbd_1375 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1375", this);
    pf_vf_mux_scbd_1376 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1376", this);
    pf_vf_mux_scbd_1377 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1377", this);
    pf_vf_mux_scbd_1378 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1378", this);
    pf_vf_mux_scbd_1379 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1379", this);
    pf_vf_mux_scbd_1380 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1380", this);
    pf_vf_mux_scbd_1381 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1381", this);
    pf_vf_mux_scbd_1382 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1382", this);
    pf_vf_mux_scbd_1383 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1383", this);
    pf_vf_mux_scbd_1384 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1384", this);
    pf_vf_mux_scbd_1385 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1385", this);
    pf_vf_mux_scbd_1386 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1386", this);
    pf_vf_mux_scbd_1387 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1387", this);
    pf_vf_mux_scbd_1388 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1388", this);
    pf_vf_mux_scbd_1389 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1389", this);
    pf_vf_mux_scbd_1390 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1390", this);
    pf_vf_mux_scbd_1391 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1391", this);
    pf_vf_mux_scbd_1392 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1392", this);
    pf_vf_mux_scbd_1393 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1393", this);
    pf_vf_mux_scbd_1394 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1394", this);
    pf_vf_mux_scbd_1395 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1395", this);
    pf_vf_mux_scbd_1396 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1396", this);
    pf_vf_mux_scbd_1397 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1397", this);
    pf_vf_mux_scbd_1398 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1398", this);
    pf_vf_mux_scbd_1399 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1399", this);
    pf_vf_mux_scbd_1400 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1400", this);
    pf_vf_mux_scbd_1401 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1401", this);
    pf_vf_mux_scbd_1402 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1402", this);
    pf_vf_mux_scbd_1403 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1403", this);
    pf_vf_mux_scbd_1404 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1404", this);
    pf_vf_mux_scbd_1405 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1405", this);
    pf_vf_mux_scbd_1406 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1406", this);
    pf_vf_mux_scbd_1407 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1407", this);
    pf_vf_mux_scbd_1408 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1408", this);
    pf_vf_mux_scbd_1409 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1409", this);
    pf_vf_mux_scbd_1410 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1410", this);
    pf_vf_mux_scbd_1411 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1411", this);
    pf_vf_mux_scbd_1412 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1412", this);
    pf_vf_mux_scbd_1413 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1413", this);
    pf_vf_mux_scbd_1414 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1414", this);
    pf_vf_mux_scbd_1415 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1415", this);
    pf_vf_mux_scbd_1416 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1416", this);
    pf_vf_mux_scbd_1417 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1417", this);
    pf_vf_mux_scbd_1418 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1418", this);
    pf_vf_mux_scbd_1419 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1419", this);
    pf_vf_mux_scbd_1420 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1420", this);
    pf_vf_mux_scbd_1421 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1421", this);
    pf_vf_mux_scbd_1422 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1422", this);
    pf_vf_mux_scbd_1423 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1423", this);
    pf_vf_mux_scbd_1424 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1424", this);
    pf_vf_mux_scbd_1425 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1425", this);
    pf_vf_mux_scbd_1426 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1426", this);
    pf_vf_mux_scbd_1427 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1427", this);
    pf_vf_mux_scbd_1428 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1428", this);
    pf_vf_mux_scbd_1429 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1429", this);
    pf_vf_mux_scbd_1430 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1430", this);
    pf_vf_mux_scbd_1431 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1431", this);
    pf_vf_mux_scbd_1432 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1432", this);
    pf_vf_mux_scbd_1433 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1433", this);
    pf_vf_mux_scbd_1434 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1434", this);
    pf_vf_mux_scbd_1435 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1435", this);
    pf_vf_mux_scbd_1436 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1436", this);
    pf_vf_mux_scbd_1437 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1437", this);
    pf_vf_mux_scbd_1438 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1438", this);
    pf_vf_mux_scbd_1439 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1439", this);
    pf_vf_mux_scbd_1440 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1440", this);
    pf_vf_mux_scbd_1441 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1441", this);
    pf_vf_mux_scbd_1442 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1442", this);
    pf_vf_mux_scbd_1443 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1443", this);
    pf_vf_mux_scbd_1444 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1444", this);
    pf_vf_mux_scbd_1445 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1445", this);
    pf_vf_mux_scbd_1446 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1446", this);
    pf_vf_mux_scbd_1447 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1447", this);
    pf_vf_mux_scbd_1448 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1448", this);
    pf_vf_mux_scbd_1449 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1449", this);
    pf_vf_mux_scbd_1450 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1450", this);
    pf_vf_mux_scbd_1451 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1451", this);
    pf_vf_mux_scbd_1452 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1452", this);
    pf_vf_mux_scbd_1453 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1453", this);
    pf_vf_mux_scbd_1454 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1454", this);
    pf_vf_mux_scbd_1455 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1455", this);
    pf_vf_mux_scbd_1456 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1456", this);
    pf_vf_mux_scbd_1457 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1457", this);
    pf_vf_mux_scbd_1458 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1458", this);
    pf_vf_mux_scbd_1459 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1459", this);
    pf_vf_mux_scbd_1460 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1460", this);
    pf_vf_mux_scbd_1461 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1461", this);
    pf_vf_mux_scbd_1462 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1462", this);
    pf_vf_mux_scbd_1463 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1463", this);
    pf_vf_mux_scbd_1464 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1464", this);
    pf_vf_mux_scbd_1465 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1465", this);
    pf_vf_mux_scbd_1466 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1466", this);
    pf_vf_mux_scbd_1467 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1467", this);
    pf_vf_mux_scbd_1468 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1468", this);
    pf_vf_mux_scbd_1469 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1469", this);
    pf_vf_mux_scbd_1470 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1470", this);
    pf_vf_mux_scbd_1471 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1471", this);
    pf_vf_mux_scbd_1472 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1472", this);
    pf_vf_mux_scbd_1473 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1473", this);
    pf_vf_mux_scbd_1474 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1474", this);
    pf_vf_mux_scbd_1475 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1475", this);
    pf_vf_mux_scbd_1476 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1476", this);
    pf_vf_mux_scbd_1477 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1477", this);
    pf_vf_mux_scbd_1478 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1478", this);
    pf_vf_mux_scbd_1479 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1479", this);
    pf_vf_mux_scbd_1480 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1480", this);
    pf_vf_mux_scbd_1481 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1481", this);
    pf_vf_mux_scbd_1482 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1482", this);
    pf_vf_mux_scbd_1483 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1483", this);
    pf_vf_mux_scbd_1484 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1484", this);
    pf_vf_mux_scbd_1485 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1485", this);
    pf_vf_mux_scbd_1486 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1486", this);
    pf_vf_mux_scbd_1487 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1487", this);
    pf_vf_mux_scbd_1488 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1488", this);
    pf_vf_mux_scbd_1489 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1489", this);
    pf_vf_mux_scbd_1490 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1490", this);
    pf_vf_mux_scbd_1491 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1491", this);
    pf_vf_mux_scbd_1492 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1492", this);
    pf_vf_mux_scbd_1493 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1493", this);
    pf_vf_mux_scbd_1494 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1494", this);
    pf_vf_mux_scbd_1495 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1495", this);
    pf_vf_mux_scbd_1496 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1496", this);
    pf_vf_mux_scbd_1497 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1497", this);
    pf_vf_mux_scbd_1498 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1498", this);
    pf_vf_mux_scbd_1499 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1499", this);
    pf_vf_mux_scbd_1500 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1500", this);
    pf_vf_mux_scbd_1501 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1501", this);
    pf_vf_mux_scbd_1502 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1502", this);
    pf_vf_mux_scbd_1503 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1503", this);
    pf_vf_mux_scbd_1504 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1504", this);
    pf_vf_mux_scbd_1505 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1505", this);
    pf_vf_mux_scbd_1506 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1506", this);
    pf_vf_mux_scbd_1507 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1507", this);
    pf_vf_mux_scbd_1508 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1508", this);
    pf_vf_mux_scbd_1509 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1509", this);
    pf_vf_mux_scbd_1510 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1510", this);
    pf_vf_mux_scbd_1511 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1511", this);
    pf_vf_mux_scbd_1512 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1512", this);
    pf_vf_mux_scbd_1513 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1513", this);
    pf_vf_mux_scbd_1514 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1514", this);
    pf_vf_mux_scbd_1515 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1515", this);
    pf_vf_mux_scbd_1516 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1516", this);
    pf_vf_mux_scbd_1517 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1517", this);
    pf_vf_mux_scbd_1518 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1518", this);
    pf_vf_mux_scbd_1519 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1519", this);
    pf_vf_mux_scbd_1520 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1520", this);
    pf_vf_mux_scbd_1521 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1521", this);
    pf_vf_mux_scbd_1522 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1522", this);
    pf_vf_mux_scbd_1523 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1523", this);
    pf_vf_mux_scbd_1524 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1524", this);
    pf_vf_mux_scbd_1525 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1525", this);
    pf_vf_mux_scbd_1526 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1526", this);
    pf_vf_mux_scbd_1527 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1527", this);
    pf_vf_mux_scbd_1528 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1528", this);
    pf_vf_mux_scbd_1529 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1529", this);
    pf_vf_mux_scbd_1530 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1530", this);
    pf_vf_mux_scbd_1531 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1531", this);
    pf_vf_mux_scbd_1532 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1532", this);
    pf_vf_mux_scbd_1533 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1533", this);
    pf_vf_mux_scbd_1534 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1534", this);
    pf_vf_mux_scbd_1535 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1535", this);
    pf_vf_mux_scbd_1536 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1536", this);
    pf_vf_mux_scbd_1537 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1537", this);
    pf_vf_mux_scbd_1538 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1538", this);
    pf_vf_mux_scbd_1539 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1539", this);
    pf_vf_mux_scbd_1540 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1540", this);
    pf_vf_mux_scbd_1541 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1541", this);
    pf_vf_mux_scbd_1542 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1542", this);
    pf_vf_mux_scbd_1543 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1543", this);
    pf_vf_mux_scbd_1544 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1544", this);
    pf_vf_mux_scbd_1545 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1545", this);
    pf_vf_mux_scbd_1546 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1546", this);
    pf_vf_mux_scbd_1547 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1547", this);
    pf_vf_mux_scbd_1548 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1548", this);
    pf_vf_mux_scbd_1549 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1549", this);
    pf_vf_mux_scbd_1550 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1550", this);
    pf_vf_mux_scbd_1551 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1551", this);
    pf_vf_mux_scbd_1552 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1552", this);
    pf_vf_mux_scbd_1553 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1553", this);
    pf_vf_mux_scbd_1554 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1554", this);
    pf_vf_mux_scbd_1555 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1555", this);
    pf_vf_mux_scbd_1556 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1556", this);
    pf_vf_mux_scbd_1557 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1557", this);
    pf_vf_mux_scbd_1558 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1558", this);
    pf_vf_mux_scbd_1559 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1559", this);
    pf_vf_mux_scbd_1560 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1560", this);
    pf_vf_mux_scbd_1561 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1561", this);
    pf_vf_mux_scbd_1562 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1562", this);
    pf_vf_mux_scbd_1563 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1563", this);
    pf_vf_mux_scbd_1564 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1564", this);
    pf_vf_mux_scbd_1565 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1565", this);
    pf_vf_mux_scbd_1566 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1566", this);
    pf_vf_mux_scbd_1567 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1567", this);
    pf_vf_mux_scbd_1568 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1568", this);
    pf_vf_mux_scbd_1569 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1569", this);
    pf_vf_mux_scbd_1570 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1570", this);
    pf_vf_mux_scbd_1571 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1571", this);
    pf_vf_mux_scbd_1572 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1572", this);
    pf_vf_mux_scbd_1573 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1573", this);
    pf_vf_mux_scbd_1574 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1574", this);
    pf_vf_mux_scbd_1575 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1575", this);
    pf_vf_mux_scbd_1576 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1576", this);
    pf_vf_mux_scbd_1577 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1577", this);
    pf_vf_mux_scbd_1578 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1578", this);
    pf_vf_mux_scbd_1579 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1579", this);
    pf_vf_mux_scbd_1580 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1580", this);
    pf_vf_mux_scbd_1581 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1581", this);
    pf_vf_mux_scbd_1582 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1582", this);
    pf_vf_mux_scbd_1583 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1583", this);
    pf_vf_mux_scbd_1584 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1584", this);
    pf_vf_mux_scbd_1585 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1585", this);
    pf_vf_mux_scbd_1586 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1586", this);
    pf_vf_mux_scbd_1587 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1587", this);
    pf_vf_mux_scbd_1588 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1588", this);
    pf_vf_mux_scbd_1589 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1589", this);
    pf_vf_mux_scbd_1590 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1590", this);
    pf_vf_mux_scbd_1591 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1591", this);
    pf_vf_mux_scbd_1592 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1592", this);
    pf_vf_mux_scbd_1593 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1593", this);
    pf_vf_mux_scbd_1594 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1594", this);
    pf_vf_mux_scbd_1595 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1595", this);
    pf_vf_mux_scbd_1596 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1596", this);
    pf_vf_mux_scbd_1597 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1597", this);
    pf_vf_mux_scbd_1598 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1598", this);
    pf_vf_mux_scbd_1599 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1599", this);
    pf_vf_mux_scbd_1600 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1600", this);
    pf_vf_mux_scbd_1601 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1601", this);
    pf_vf_mux_scbd_1602 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1602", this);
    pf_vf_mux_scbd_1603 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1603", this);
    pf_vf_mux_scbd_1604 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1604", this);
    pf_vf_mux_scbd_1605 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1605", this);
    pf_vf_mux_scbd_1606 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1606", this);
    pf_vf_mux_scbd_1607 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1607", this);
    pf_vf_mux_scbd_1608 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1608", this);
    pf_vf_mux_scbd_1609 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1609", this);
    pf_vf_mux_scbd_1610 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1610", this);
    pf_vf_mux_scbd_1611 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1611", this);
    pf_vf_mux_scbd_1612 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1612", this);
    pf_vf_mux_scbd_1613 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1613", this);
    pf_vf_mux_scbd_1614 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1614", this);
    pf_vf_mux_scbd_1615 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1615", this);
    pf_vf_mux_scbd_1616 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1616", this);
    pf_vf_mux_scbd_1617 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1617", this);
    pf_vf_mux_scbd_1618 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1618", this);
    pf_vf_mux_scbd_1619 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1619", this);
    pf_vf_mux_scbd_1620 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1620", this);
    pf_vf_mux_scbd_1621 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1621", this);
    pf_vf_mux_scbd_1622 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1622", this);
    pf_vf_mux_scbd_1623 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1623", this);
    pf_vf_mux_scbd_1624 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1624", this);
    pf_vf_mux_scbd_1625 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1625", this);
    pf_vf_mux_scbd_1626 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1626", this);
    pf_vf_mux_scbd_1627 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1627", this);
    pf_vf_mux_scbd_1628 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1628", this);
    pf_vf_mux_scbd_1629 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1629", this);
    pf_vf_mux_scbd_1630 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1630", this);
    pf_vf_mux_scbd_1631 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1631", this);
    pf_vf_mux_scbd_1632 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1632", this);
    pf_vf_mux_scbd_1633 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1633", this);
    pf_vf_mux_scbd_1634 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1634", this);
    pf_vf_mux_scbd_1635 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1635", this);
    pf_vf_mux_scbd_1636 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1636", this);
    pf_vf_mux_scbd_1637 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1637", this);
    pf_vf_mux_scbd_1638 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1638", this);
    pf_vf_mux_scbd_1639 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1639", this);
    pf_vf_mux_scbd_1640 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1640", this);
    pf_vf_mux_scbd_1641 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1641", this);
    pf_vf_mux_scbd_1642 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1642", this);
    pf_vf_mux_scbd_1643 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1643", this);
    pf_vf_mux_scbd_1644 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1644", this);
    pf_vf_mux_scbd_1645 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1645", this);
    pf_vf_mux_scbd_1646 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1646", this);
    pf_vf_mux_scbd_1647 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1647", this);
    pf_vf_mux_scbd_1648 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1648", this);
    pf_vf_mux_scbd_1649 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1649", this);
    pf_vf_mux_scbd_1650 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1650", this);
    pf_vf_mux_scbd_1651 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1651", this);
    pf_vf_mux_scbd_1652 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1652", this);
    pf_vf_mux_scbd_1653 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1653", this);
    pf_vf_mux_scbd_1654 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1654", this);
    pf_vf_mux_scbd_1655 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1655", this);
    pf_vf_mux_scbd_1656 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1656", this);
    pf_vf_mux_scbd_1657 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1657", this);
    pf_vf_mux_scbd_1658 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1658", this);
    pf_vf_mux_scbd_1659 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1659", this);
    pf_vf_mux_scbd_1660 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1660", this);
    pf_vf_mux_scbd_1661 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1661", this);
    pf_vf_mux_scbd_1662 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1662", this);
    pf_vf_mux_scbd_1663 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1663", this);
    pf_vf_mux_scbd_1664 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1664", this);
    pf_vf_mux_scbd_1665 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1665", this);
    pf_vf_mux_scbd_1666 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1666", this);
    pf_vf_mux_scbd_1667 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1667", this);
    pf_vf_mux_scbd_1668 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1668", this);
    pf_vf_mux_scbd_1669 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1669", this);
    pf_vf_mux_scbd_1670 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1670", this);
    pf_vf_mux_scbd_1671 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1671", this);
    pf_vf_mux_scbd_1672 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1672", this);
    pf_vf_mux_scbd_1673 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1673", this);
    pf_vf_mux_scbd_1674 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1674", this);
    pf_vf_mux_scbd_1675 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1675", this);
    pf_vf_mux_scbd_1676 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1676", this);
    pf_vf_mux_scbd_1677 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1677", this);
    pf_vf_mux_scbd_1678 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1678", this);
    pf_vf_mux_scbd_1679 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1679", this);
    pf_vf_mux_scbd_1680 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1680", this);
    pf_vf_mux_scbd_1681 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1681", this);
    pf_vf_mux_scbd_1682 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1682", this);
    pf_vf_mux_scbd_1683 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1683", this);
    pf_vf_mux_scbd_1684 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1684", this);
    pf_vf_mux_scbd_1685 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1685", this);
    pf_vf_mux_scbd_1686 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1686", this);
    pf_vf_mux_scbd_1687 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1687", this);
    pf_vf_mux_scbd_1688 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1688", this);
    pf_vf_mux_scbd_1689 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1689", this);
    pf_vf_mux_scbd_1690 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1690", this);
    pf_vf_mux_scbd_1691 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1691", this);
    pf_vf_mux_scbd_1692 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1692", this);
    pf_vf_mux_scbd_1693 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1693", this);
    pf_vf_mux_scbd_1694 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1694", this);
    pf_vf_mux_scbd_1695 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1695", this);
    pf_vf_mux_scbd_1696 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1696", this);
    pf_vf_mux_scbd_1697 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1697", this);
    pf_vf_mux_scbd_1698 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1698", this);
    pf_vf_mux_scbd_1699 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1699", this);
    pf_vf_mux_scbd_1700 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1700", this);
    pf_vf_mux_scbd_1701 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1701", this);
    pf_vf_mux_scbd_1702 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1702", this);
    pf_vf_mux_scbd_1703 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1703", this);
    pf_vf_mux_scbd_1704 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1704", this);
    pf_vf_mux_scbd_1705 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1705", this);
    pf_vf_mux_scbd_1706 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1706", this);
    pf_vf_mux_scbd_1707 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1707", this);
    pf_vf_mux_scbd_1708 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1708", this);
    pf_vf_mux_scbd_1709 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1709", this);
    pf_vf_mux_scbd_1710 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1710", this);
    pf_vf_mux_scbd_1711 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1711", this);
    pf_vf_mux_scbd_1712 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1712", this);
    pf_vf_mux_scbd_1713 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1713", this);
    pf_vf_mux_scbd_1714 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1714", this);
    pf_vf_mux_scbd_1715 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1715", this);
    pf_vf_mux_scbd_1716 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1716", this);
    pf_vf_mux_scbd_1717 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1717", this);
    pf_vf_mux_scbd_1718 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1718", this);
    pf_vf_mux_scbd_1719 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1719", this);
    pf_vf_mux_scbd_1720 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1720", this);
    pf_vf_mux_scbd_1721 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1721", this);
    pf_vf_mux_scbd_1722 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1722", this);
    pf_vf_mux_scbd_1723 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1723", this);
    pf_vf_mux_scbd_1724 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1724", this);
    pf_vf_mux_scbd_1725 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1725", this);
    pf_vf_mux_scbd_1726 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1726", this);
    pf_vf_mux_scbd_1727 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1727", this);
    pf_vf_mux_scbd_1728 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1728", this);
    pf_vf_mux_scbd_1729 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1729", this);
    pf_vf_mux_scbd_1730 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1730", this);
    pf_vf_mux_scbd_1731 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1731", this);
    pf_vf_mux_scbd_1732 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1732", this);
    pf_vf_mux_scbd_1733 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1733", this);
    pf_vf_mux_scbd_1734 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1734", this);
    pf_vf_mux_scbd_1735 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1735", this);
    pf_vf_mux_scbd_1736 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1736", this);
    pf_vf_mux_scbd_1737 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1737", this);
    pf_vf_mux_scbd_1738 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1738", this);
    pf_vf_mux_scbd_1739 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1739", this);
    pf_vf_mux_scbd_1740 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1740", this);
    pf_vf_mux_scbd_1741 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1741", this);
    pf_vf_mux_scbd_1742 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1742", this);
    pf_vf_mux_scbd_1743 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1743", this);
    pf_vf_mux_scbd_1744 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1744", this);
    pf_vf_mux_scbd_1745 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1745", this);
    pf_vf_mux_scbd_1746 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1746", this);
    pf_vf_mux_scbd_1747 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1747", this);
    pf_vf_mux_scbd_1748 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1748", this);
    pf_vf_mux_scbd_1749 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1749", this);
    pf_vf_mux_scbd_1750 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1750", this);
    pf_vf_mux_scbd_1751 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1751", this);
    pf_vf_mux_scbd_1752 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1752", this);
    pf_vf_mux_scbd_1753 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1753", this);
    pf_vf_mux_scbd_1754 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1754", this);
    pf_vf_mux_scbd_1755 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1755", this);
    pf_vf_mux_scbd_1756 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1756", this);
    pf_vf_mux_scbd_1757 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1757", this);
    pf_vf_mux_scbd_1758 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1758", this);
    pf_vf_mux_scbd_1759 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1759", this);
    pf_vf_mux_scbd_1760 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1760", this);
    pf_vf_mux_scbd_1761 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1761", this);
    pf_vf_mux_scbd_1762 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1762", this);
    pf_vf_mux_scbd_1763 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1763", this);
    pf_vf_mux_scbd_1764 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1764", this);
    pf_vf_mux_scbd_1765 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1765", this);
    pf_vf_mux_scbd_1766 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1766", this);
    pf_vf_mux_scbd_1767 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1767", this);
    pf_vf_mux_scbd_1768 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1768", this);
    pf_vf_mux_scbd_1769 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1769", this);
    pf_vf_mux_scbd_1770 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1770", this);
    pf_vf_mux_scbd_1771 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1771", this);
    pf_vf_mux_scbd_1772 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1772", this);
    pf_vf_mux_scbd_1773 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1773", this);
    pf_vf_mux_scbd_1774 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1774", this);
    pf_vf_mux_scbd_1775 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1775", this);
    pf_vf_mux_scbd_1776 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1776", this);
    pf_vf_mux_scbd_1777 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1777", this);
    pf_vf_mux_scbd_1778 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1778", this);
    pf_vf_mux_scbd_1779 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1779", this);
    pf_vf_mux_scbd_1780 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1780", this);
    pf_vf_mux_scbd_1781 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1781", this);
    pf_vf_mux_scbd_1782 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1782", this);
    pf_vf_mux_scbd_1783 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1783", this);
    pf_vf_mux_scbd_1784 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1784", this);
    pf_vf_mux_scbd_1785 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1785", this);
    pf_vf_mux_scbd_1786 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1786", this);
    pf_vf_mux_scbd_1787 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1787", this);
    pf_vf_mux_scbd_1788 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1788", this);
    pf_vf_mux_scbd_1789 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1789", this);
    pf_vf_mux_scbd_1790 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1790", this);
    pf_vf_mux_scbd_1791 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1791", this);
    pf_vf_mux_scbd_1792 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1792", this);
    pf_vf_mux_scbd_1793 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1793", this);
    pf_vf_mux_scbd_1794 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1794", this);
    pf_vf_mux_scbd_1795 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1795", this);
    pf_vf_mux_scbd_1796 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1796", this);
    pf_vf_mux_scbd_1797 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1797", this);
    pf_vf_mux_scbd_1798 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1798", this);
    pf_vf_mux_scbd_1799 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1799", this);
    pf_vf_mux_scbd_1800 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1800", this);
    pf_vf_mux_scbd_1801 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1801", this);
    pf_vf_mux_scbd_1802 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1802", this);
    pf_vf_mux_scbd_1803 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1803", this);
    pf_vf_mux_scbd_1804 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1804", this);
    pf_vf_mux_scbd_1805 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1805", this);
    pf_vf_mux_scbd_1806 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1806", this);
    pf_vf_mux_scbd_1807 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1807", this);
    pf_vf_mux_scbd_1808 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1808", this);
    pf_vf_mux_scbd_1809 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1809", this);
    pf_vf_mux_scbd_1810 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1810", this);
    pf_vf_mux_scbd_1811 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1811", this);
    pf_vf_mux_scbd_1812 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1812", this);
    pf_vf_mux_scbd_1813 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1813", this);
    pf_vf_mux_scbd_1814 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1814", this);
    pf_vf_mux_scbd_1815 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1815", this);
    pf_vf_mux_scbd_1816 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1816", this);
    pf_vf_mux_scbd_1817 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1817", this);
    pf_vf_mux_scbd_1818 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1818", this);
    pf_vf_mux_scbd_1819 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1819", this);
    pf_vf_mux_scbd_1820 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1820", this);
    pf_vf_mux_scbd_1821 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1821", this);
    pf_vf_mux_scbd_1822 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1822", this);
    pf_vf_mux_scbd_1823 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1823", this);
    pf_vf_mux_scbd_1824 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1824", this);
    pf_vf_mux_scbd_1825 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1825", this);
    pf_vf_mux_scbd_1826 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1826", this);
    pf_vf_mux_scbd_1827 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1827", this);
    pf_vf_mux_scbd_1828 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1828", this);
    pf_vf_mux_scbd_1829 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1829", this);
    pf_vf_mux_scbd_1830 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1830", this);
    pf_vf_mux_scbd_1831 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1831", this);
    pf_vf_mux_scbd_1832 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1832", this);
    pf_vf_mux_scbd_1833 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1833", this);
    pf_vf_mux_scbd_1834 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1834", this);
    pf_vf_mux_scbd_1835 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1835", this);
    pf_vf_mux_scbd_1836 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1836", this);
    pf_vf_mux_scbd_1837 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1837", this);
    pf_vf_mux_scbd_1838 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1838", this);
    pf_vf_mux_scbd_1839 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1839", this);
    pf_vf_mux_scbd_1840 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1840", this);
    pf_vf_mux_scbd_1841 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1841", this);
    pf_vf_mux_scbd_1842 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1842", this);
    pf_vf_mux_scbd_1843 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1843", this);
    pf_vf_mux_scbd_1844 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1844", this);
    pf_vf_mux_scbd_1845 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1845", this);
    pf_vf_mux_scbd_1846 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1846", this);
    pf_vf_mux_scbd_1847 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1847", this);
    pf_vf_mux_scbd_1848 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1848", this);
    pf_vf_mux_scbd_1849 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1849", this);
    pf_vf_mux_scbd_1850 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1850", this);
    pf_vf_mux_scbd_1851 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1851", this);
    pf_vf_mux_scbd_1852 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1852", this);
    pf_vf_mux_scbd_1853 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1853", this);
    pf_vf_mux_scbd_1854 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1854", this);
    pf_vf_mux_scbd_1855 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1855", this);
    pf_vf_mux_scbd_1856 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1856", this);
    pf_vf_mux_scbd_1857 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1857", this);
    pf_vf_mux_scbd_1858 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1858", this);
    pf_vf_mux_scbd_1859 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1859", this);
    pf_vf_mux_scbd_1860 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1860", this);
    pf_vf_mux_scbd_1861 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1861", this);
    pf_vf_mux_scbd_1862 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1862", this);
    pf_vf_mux_scbd_1863 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1863", this);
    pf_vf_mux_scbd_1864 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1864", this);
    pf_vf_mux_scbd_1865 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1865", this);
    pf_vf_mux_scbd_1866 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1866", this);
    pf_vf_mux_scbd_1867 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1867", this);
    pf_vf_mux_scbd_1868 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1868", this);
    pf_vf_mux_scbd_1869 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1869", this);
    pf_vf_mux_scbd_1870 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1870", this);
    pf_vf_mux_scbd_1871 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1871", this);
    pf_vf_mux_scbd_1872 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1872", this);
    pf_vf_mux_scbd_1873 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1873", this);
    pf_vf_mux_scbd_1874 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1874", this);
    pf_vf_mux_scbd_1875 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1875", this);
    pf_vf_mux_scbd_1876 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1876", this);
    pf_vf_mux_scbd_1877 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1877", this);
    pf_vf_mux_scbd_1878 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1878", this);
    pf_vf_mux_scbd_1879 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1879", this);
    pf_vf_mux_scbd_1880 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1880", this);
    pf_vf_mux_scbd_1881 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1881", this);
    pf_vf_mux_scbd_1882 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1882", this);
    pf_vf_mux_scbd_1883 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1883", this);
    pf_vf_mux_scbd_1884 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1884", this);
    pf_vf_mux_scbd_1885 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1885", this);
    pf_vf_mux_scbd_1886 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1886", this);
    pf_vf_mux_scbd_1887 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1887", this);
    pf_vf_mux_scbd_1888 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1888", this);
    pf_vf_mux_scbd_1889 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1889", this);
    pf_vf_mux_scbd_1890 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1890", this);
    pf_vf_mux_scbd_1891 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1891", this);
    pf_vf_mux_scbd_1892 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1892", this);
    pf_vf_mux_scbd_1893 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1893", this);
    pf_vf_mux_scbd_1894 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1894", this);
    pf_vf_mux_scbd_1895 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1895", this);
    pf_vf_mux_scbd_1896 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1896", this);
    pf_vf_mux_scbd_1897 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1897", this);
    pf_vf_mux_scbd_1898 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1898", this);
    pf_vf_mux_scbd_1899 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1899", this);
    pf_vf_mux_scbd_1900 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1900", this);
    pf_vf_mux_scbd_1901 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1901", this);
    pf_vf_mux_scbd_1902 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1902", this);
    pf_vf_mux_scbd_1903 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1903", this);
    pf_vf_mux_scbd_1904 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1904", this);
    pf_vf_mux_scbd_1905 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1905", this);
    pf_vf_mux_scbd_1906 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1906", this);
    pf_vf_mux_scbd_1907 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1907", this);
    pf_vf_mux_scbd_1908 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1908", this);
    pf_vf_mux_scbd_1909 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1909", this);
    pf_vf_mux_scbd_1910 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1910", this);
    pf_vf_mux_scbd_1911 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1911", this);
    pf_vf_mux_scbd_1912 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1912", this);
    pf_vf_mux_scbd_1913 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1913", this);
    pf_vf_mux_scbd_1914 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1914", this);
    pf_vf_mux_scbd_1915 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1915", this);
    pf_vf_mux_scbd_1916 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1916", this);
    pf_vf_mux_scbd_1917 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1917", this);
    pf_vf_mux_scbd_1918 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1918", this);
    pf_vf_mux_scbd_1919 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1919", this);
    pf_vf_mux_scbd_1920 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1920", this);
    pf_vf_mux_scbd_1921 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1921", this);
    pf_vf_mux_scbd_1922 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1922", this);
    pf_vf_mux_scbd_1923 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1923", this);
    pf_vf_mux_scbd_1924 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1924", this);
    pf_vf_mux_scbd_1925 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1925", this);
    pf_vf_mux_scbd_1926 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1926", this);
    pf_vf_mux_scbd_1927 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1927", this);
    pf_vf_mux_scbd_1928 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1928", this);
    pf_vf_mux_scbd_1929 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1929", this);
    pf_vf_mux_scbd_1930 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1930", this);
    pf_vf_mux_scbd_1931 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1931", this);
    pf_vf_mux_scbd_1932 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1932", this);
    pf_vf_mux_scbd_1933 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1933", this);
    pf_vf_mux_scbd_1934 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1934", this);
    pf_vf_mux_scbd_1935 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1935", this);
    pf_vf_mux_scbd_1936 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1936", this);
    pf_vf_mux_scbd_1937 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1937", this);
    pf_vf_mux_scbd_1938 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1938", this);
    pf_vf_mux_scbd_1939 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1939", this);
    pf_vf_mux_scbd_1940 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1940", this);
    pf_vf_mux_scbd_1941 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1941", this);
    pf_vf_mux_scbd_1942 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1942", this);
    pf_vf_mux_scbd_1943 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1943", this);
    pf_vf_mux_scbd_1944 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1944", this);
    pf_vf_mux_scbd_1945 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1945", this);
    pf_vf_mux_scbd_1946 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1946", this);
    pf_vf_mux_scbd_1947 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1947", this);
    pf_vf_mux_scbd_1948 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1948", this);
    pf_vf_mux_scbd_1949 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1949", this);
    pf_vf_mux_scbd_1950 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1950", this);
    pf_vf_mux_scbd_1951 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1951", this);
    pf_vf_mux_scbd_1952 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1952", this);
    pf_vf_mux_scbd_1953 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1953", this);
    pf_vf_mux_scbd_1954 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1954", this);
    pf_vf_mux_scbd_1955 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1955", this);
    pf_vf_mux_scbd_1956 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1956", this);
    pf_vf_mux_scbd_1957 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1957", this);
    pf_vf_mux_scbd_1958 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1958", this);
    pf_vf_mux_scbd_1959 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1959", this);
    pf_vf_mux_scbd_1960 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1960", this);
    pf_vf_mux_scbd_1961 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1961", this);
    pf_vf_mux_scbd_1962 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1962", this);
    pf_vf_mux_scbd_1963 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1963", this);
    pf_vf_mux_scbd_1964 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1964", this);
    pf_vf_mux_scbd_1965 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1965", this);
    pf_vf_mux_scbd_1966 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1966", this);
    pf_vf_mux_scbd_1967 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1967", this);
    pf_vf_mux_scbd_1968 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1968", this);
    pf_vf_mux_scbd_1969 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1969", this);
    pf_vf_mux_scbd_1970 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1970", this);
    pf_vf_mux_scbd_1971 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1971", this);
    pf_vf_mux_scbd_1972 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1972", this);
    pf_vf_mux_scbd_1973 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1973", this);
    pf_vf_mux_scbd_1974 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1974", this);
    pf_vf_mux_scbd_1975 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1975", this);
    pf_vf_mux_scbd_1976 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1976", this);
    pf_vf_mux_scbd_1977 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1977", this);
    pf_vf_mux_scbd_1978 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1978", this);
    pf_vf_mux_scbd_1979 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1979", this);
    pf_vf_mux_scbd_1980 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1980", this);
    pf_vf_mux_scbd_1981 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1981", this);
    pf_vf_mux_scbd_1982 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1982", this);
    pf_vf_mux_scbd_1983 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1983", this);
    pf_vf_mux_scbd_1984 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1984", this);
    pf_vf_mux_scbd_1985 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1985", this);
    pf_vf_mux_scbd_1986 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1986", this);
    pf_vf_mux_scbd_1987 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1987", this);
    pf_vf_mux_scbd_1988 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1988", this);
    pf_vf_mux_scbd_1989 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1989", this);
    pf_vf_mux_scbd_1990 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1990", this);
    pf_vf_mux_scbd_1991 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1991", this);
    pf_vf_mux_scbd_1992 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1992", this);
    pf_vf_mux_scbd_1993 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1993", this);
    pf_vf_mux_scbd_1994 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1994", this);
    pf_vf_mux_scbd_1995 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1995", this);
    pf_vf_mux_scbd_1996 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1996", this);
    pf_vf_mux_scbd_1997 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1997", this);
    pf_vf_mux_scbd_1998 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1998", this);
    pf_vf_mux_scbd_1999 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1999", this);
    pf_vf_mux_scbd_2000 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2000", this);
    pf_vf_mux_scbd_2001 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2001", this);
    pf_vf_mux_scbd_2002 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2002", this);
    pf_vf_mux_scbd_2003 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2003", this);
    pf_vf_mux_scbd_2004 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2004", this);
    pf_vf_mux_scbd_2005 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2005", this);
    pf_vf_mux_scbd_2006 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2006", this);
    pf_vf_mux_scbd_2007 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2007", this);
    pf_vf_mux_scbd_2008 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2008", this);
    pf_vf_mux_scbd_2009 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2009", this);
    pf_vf_mux_scbd_2010 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2010", this);
    pf_vf_mux_scbd_2011 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2011", this);
    pf_vf_mux_scbd_2012 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2012", this);
    pf_vf_mux_scbd_2013 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2013", this);
    pf_vf_mux_scbd_2014 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2014", this);
    pf_vf_mux_scbd_2015 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2015", this);
    pf_vf_mux_scbd_2016 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2016", this);
    pf_vf_mux_scbd_2017 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2017", this);
    pf_vf_mux_scbd_2018 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2018", this);
    pf_vf_mux_scbd_2019 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2019", this);
    pf_vf_mux_scbd_2020 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2020", this);
    pf_vf_mux_scbd_2021 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2021", this);
    pf_vf_mux_scbd_2022 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2022", this);
    pf_vf_mux_scbd_2023 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2023", this);
    pf_vf_mux_scbd_2024 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2024", this);
    pf_vf_mux_scbd_2025 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2025", this);
    pf_vf_mux_scbd_2026 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2026", this);
    pf_vf_mux_scbd_2027 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2027", this);
    pf_vf_mux_scbd_2028 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2028", this);
    pf_vf_mux_scbd_2029 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2029", this);
    pf_vf_mux_scbd_2030 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2030", this);
    pf_vf_mux_scbd_2031 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2031", this);
    pf_vf_mux_scbd_2032 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2032", this);
    pf_vf_mux_scbd_2033 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2033", this);
    pf_vf_mux_scbd_2034 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2034", this);
    pf_vf_mux_scbd_2035 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2035", this);
    pf_vf_mux_scbd_2036 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2036", this);
    pf_vf_mux_scbd_2037 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2037", this);
    pf_vf_mux_scbd_2038 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2038", this);
    pf_vf_mux_scbd_2039 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2039", this);
    pf_vf_mux_scbd_2040 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2040", this);
    pf_vf_mux_scbd_2041 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2041", this);
    pf_vf_mux_scbd_2042 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2042", this);
    pf_vf_mux_scbd_2043 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2043", this);
    pf_vf_mux_scbd_2044 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2044", this);
    pf_vf_mux_scbd_2045 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2045", this);
    pf_vf_mux_scbd_2046 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2046", this);
    pf_vf_mux_scbd_2047 = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2047", this);
    `endif
    pf_vf_mux_scbd_0_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_0_up", this);
    pf_vf_mux_scbd_1_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1_up", this);
    pf_vf_mux_scbd_2_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2_up", this);
    pf_vf_mux_scbd_3_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_3_up", this);
    pf_vf_mux_scbd_4_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_4_up", this);
    pf_vf_mux_scbd_5_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_5_up", this);
    pf_vf_mux_scbd_6_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_6_up", this);
    pf_vf_mux_scbd_7_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_7_up", this);
    pf_vf_mux_scbd_8_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_8_up", this);
    pf_vf_mux_scbd_9_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_9_up", this);
    pf_vf_mux_scbd_10_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_10_up", this);
    pf_vf_mux_scbd_11_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_11_up", this);
    pf_vf_mux_scbd_12_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_12_up", this);
    pf_vf_mux_scbd_13_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_13_up", this);
    pf_vf_mux_scbd_14_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_14_up", this);
    pf_vf_mux_scbd_15_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_15_up", this);
     `ifdef TB_CONFIG_2
    pf_vf_mux_scbd_16_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_16_up", this);
    pf_vf_mux_scbd_17_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_17_up", this);
    pf_vf_mux_scbd_18_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_18_up", this);
    pf_vf_mux_scbd_19_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_19_up", this);
    pf_vf_mux_scbd_20_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_20_up", this);
    pf_vf_mux_scbd_21_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_21_up", this);
    pf_vf_mux_scbd_22_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_22_up", this);
    pf_vf_mux_scbd_23_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_23_up", this);
     `elsif TB_CONFIG_3
    pf_vf_mux_scbd_16_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_16_up", this);
    pf_vf_mux_scbd_17_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_17_up", this);
    pf_vf_mux_scbd_18_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_18_up", this);
    pf_vf_mux_scbd_19_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_19_up", this);
    pf_vf_mux_scbd_20_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_20_up", this);
    pf_vf_mux_scbd_21_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_21_up", this);
    pf_vf_mux_scbd_22_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_22_up", this);
    pf_vf_mux_scbd_23_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_23_up", this);
    pf_vf_mux_scbd_24_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_24_up", this);
    pf_vf_mux_scbd_25_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_25_up", this);
    pf_vf_mux_scbd_26_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_26_up", this);
    pf_vf_mux_scbd_27_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_27_up", this);
    pf_vf_mux_scbd_28_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_28_up", this);
    pf_vf_mux_scbd_29_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_29_up", this);
    pf_vf_mux_scbd_30_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_30_up", this);
    pf_vf_mux_scbd_31_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_31_up", this);
    `elsif TB_CONFIG_4
    pf_vf_mux_scbd_16_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_16_up", this);
    pf_vf_mux_scbd_17_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_17_up", this);
    pf_vf_mux_scbd_18_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_18_up", this);
    pf_vf_mux_scbd_19_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_19_up", this);
    pf_vf_mux_scbd_20_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_20_up", this);
    pf_vf_mux_scbd_21_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_21_up", this);
    pf_vf_mux_scbd_22_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_22_up", this);
    pf_vf_mux_scbd_23_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_23_up", this);
    pf_vf_mux_scbd_24_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_24_up", this);
    pf_vf_mux_scbd_25_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_25_up", this);
    pf_vf_mux_scbd_26_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_26_up", this);
    pf_vf_mux_scbd_27_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_27_up", this);
    pf_vf_mux_scbd_28_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_28_up", this);
    pf_vf_mux_scbd_29_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_29_up", this);
    pf_vf_mux_scbd_30_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_30_up", this);
    pf_vf_mux_scbd_31_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_31_up", this);
    pf_vf_mux_scbd_32_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_32_up", this);
    pf_vf_mux_scbd_33_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_33_up", this);
    pf_vf_mux_scbd_34_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_34_up", this);
    pf_vf_mux_scbd_35_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_35_up", this);
    pf_vf_mux_scbd_36_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_36_up", this);
    pf_vf_mux_scbd_37_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_37_up", this);
    pf_vf_mux_scbd_38_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_38_up", this);
    pf_vf_mux_scbd_39_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_39_up", this);
    pf_vf_mux_scbd_40_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_40_up", this);
    pf_vf_mux_scbd_41_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_41_up", this);
    pf_vf_mux_scbd_42_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_42_up", this);
    pf_vf_mux_scbd_43_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_43_up", this);
    pf_vf_mux_scbd_44_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_44_up", this);
    pf_vf_mux_scbd_45_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_45_up", this);
    pf_vf_mux_scbd_46_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_46_up", this);
    pf_vf_mux_scbd_47_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_47_up", this);
    pf_vf_mux_scbd_48_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_48_up", this);
    pf_vf_mux_scbd_49_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_49_up", this);
    pf_vf_mux_scbd_50_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_50_up", this);
    pf_vf_mux_scbd_51_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_51_up", this);
    pf_vf_mux_scbd_52_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_52_up", this);
    pf_vf_mux_scbd_53_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_53_up", this);
    pf_vf_mux_scbd_54_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_54_up", this);
    pf_vf_mux_scbd_55_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_55_up", this);
    pf_vf_mux_scbd_56_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_56_up", this);
    pf_vf_mux_scbd_57_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_57_up", this);
    pf_vf_mux_scbd_58_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_58_up", this);
    pf_vf_mux_scbd_59_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_59_up", this);
    pf_vf_mux_scbd_60_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_60_up", this);
    pf_vf_mux_scbd_61_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_61_up", this);
    pf_vf_mux_scbd_62_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_62_up", this);
    pf_vf_mux_scbd_63_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_63_up", this);
    pf_vf_mux_scbd_64_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_64_up", this);
    pf_vf_mux_scbd_65_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_65_up", this);
    pf_vf_mux_scbd_66_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_66_up", this);
    pf_vf_mux_scbd_67_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_67_up", this);
    pf_vf_mux_scbd_68_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_68_up", this);
    pf_vf_mux_scbd_69_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_69_up", this);
    pf_vf_mux_scbd_70_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_70_up", this);
    pf_vf_mux_scbd_71_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_71_up", this);
    pf_vf_mux_scbd_72_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_72_up", this);
    pf_vf_mux_scbd_73_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_73_up", this);
    pf_vf_mux_scbd_74_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_74_up", this);
    pf_vf_mux_scbd_75_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_75_up", this);
    pf_vf_mux_scbd_76_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_76_up", this);
    pf_vf_mux_scbd_77_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_77_up", this);
    pf_vf_mux_scbd_78_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_78_up", this);
    pf_vf_mux_scbd_79_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_79_up", this);
    pf_vf_mux_scbd_80_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_80_up", this);
    pf_vf_mux_scbd_81_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_81_up", this);
    pf_vf_mux_scbd_82_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_82_up", this);
    pf_vf_mux_scbd_83_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_83_up", this);
    pf_vf_mux_scbd_84_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_84_up", this);
    pf_vf_mux_scbd_85_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_85_up", this);
    pf_vf_mux_scbd_86_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_86_up", this);
    pf_vf_mux_scbd_87_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_87_up", this);
    pf_vf_mux_scbd_88_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_88_up", this);
    pf_vf_mux_scbd_89_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_89_up", this);
    pf_vf_mux_scbd_90_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_90_up", this);
    pf_vf_mux_scbd_91_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_91_up", this);
    pf_vf_mux_scbd_92_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_92_up", this);
    pf_vf_mux_scbd_93_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_93_up", this);
    pf_vf_mux_scbd_94_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_94_up", this);
    pf_vf_mux_scbd_95_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_95_up", this);
    pf_vf_mux_scbd_96_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_96_up", this);
    pf_vf_mux_scbd_97_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_97_up", this);
    pf_vf_mux_scbd_98_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_98_up", this);
    pf_vf_mux_scbd_99_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_99_up", this);
    pf_vf_mux_scbd_100_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_100_up", this);
    pf_vf_mux_scbd_101_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_101_up", this);
    pf_vf_mux_scbd_102_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_102_up", this);
    pf_vf_mux_scbd_103_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_103_up", this);
    pf_vf_mux_scbd_104_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_104_up", this);
    pf_vf_mux_scbd_105_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_105_up", this);
    pf_vf_mux_scbd_106_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_106_up", this);
    pf_vf_mux_scbd_107_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_107_up", this);
    pf_vf_mux_scbd_108_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_108_up", this);
    pf_vf_mux_scbd_109_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_109_up", this);
    pf_vf_mux_scbd_110_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_110_up", this);
    pf_vf_mux_scbd_111_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_111_up", this);
    pf_vf_mux_scbd_112_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_112_up", this);
    pf_vf_mux_scbd_113_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_113_up", this);
    pf_vf_mux_scbd_114_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_114_up", this);
    pf_vf_mux_scbd_115_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_115_up", this);
    pf_vf_mux_scbd_116_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_116_up", this);
    pf_vf_mux_scbd_117_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_117_up", this);
    pf_vf_mux_scbd_118_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_118_up", this);
    pf_vf_mux_scbd_119_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_119_up", this);
    pf_vf_mux_scbd_120_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_120_up", this);
    pf_vf_mux_scbd_121_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_121_up", this);
    pf_vf_mux_scbd_122_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_122_up", this);
    pf_vf_mux_scbd_123_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_123_up", this);
    pf_vf_mux_scbd_124_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_124_up", this);
    pf_vf_mux_scbd_125_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_125_up", this);
    pf_vf_mux_scbd_126_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_126_up", this);
    pf_vf_mux_scbd_127_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_127_up", this);
    pf_vf_mux_scbd_128_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_128_up", this);
    pf_vf_mux_scbd_129_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_129_up", this);
    pf_vf_mux_scbd_130_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_130_up", this);
    pf_vf_mux_scbd_131_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_131_up", this);
    pf_vf_mux_scbd_132_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_132_up", this);
    pf_vf_mux_scbd_133_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_133_up", this);
    pf_vf_mux_scbd_134_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_134_up", this);
    pf_vf_mux_scbd_135_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_135_up", this);
    pf_vf_mux_scbd_136_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_136_up", this);
    pf_vf_mux_scbd_137_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_137_up", this);
    pf_vf_mux_scbd_138_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_138_up", this);
    pf_vf_mux_scbd_139_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_139_up", this);
    pf_vf_mux_scbd_140_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_140_up", this);
    pf_vf_mux_scbd_141_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_141_up", this);
    pf_vf_mux_scbd_142_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_142_up", this);
    pf_vf_mux_scbd_143_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_143_up", this);
    pf_vf_mux_scbd_144_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_144_up", this);
    pf_vf_mux_scbd_145_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_145_up", this);
    pf_vf_mux_scbd_146_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_146_up", this);
    pf_vf_mux_scbd_147_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_147_up", this);
    pf_vf_mux_scbd_148_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_148_up", this);
    pf_vf_mux_scbd_149_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_149_up", this);
    pf_vf_mux_scbd_150_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_150_up", this);
    pf_vf_mux_scbd_151_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_151_up", this);
    pf_vf_mux_scbd_152_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_152_up", this);
    pf_vf_mux_scbd_153_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_153_up", this);
    pf_vf_mux_scbd_154_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_154_up", this);
    pf_vf_mux_scbd_155_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_155_up", this);
    pf_vf_mux_scbd_156_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_156_up", this);
    pf_vf_mux_scbd_157_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_157_up", this);
    pf_vf_mux_scbd_158_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_158_up", this);
    pf_vf_mux_scbd_159_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_159_up", this);
    pf_vf_mux_scbd_160_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_160_up", this);
    pf_vf_mux_scbd_161_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_161_up", this);
    pf_vf_mux_scbd_162_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_162_up", this);
    pf_vf_mux_scbd_163_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_163_up", this);
    pf_vf_mux_scbd_164_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_164_up", this);
    pf_vf_mux_scbd_165_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_165_up", this);
    pf_vf_mux_scbd_166_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_166_up", this);
    pf_vf_mux_scbd_167_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_167_up", this);
    pf_vf_mux_scbd_168_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_168_up", this);
    pf_vf_mux_scbd_169_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_169_up", this);
    pf_vf_mux_scbd_170_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_170_up", this);
    pf_vf_mux_scbd_171_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_171_up", this);
    pf_vf_mux_scbd_172_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_172_up", this);
    pf_vf_mux_scbd_173_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_173_up", this);
    pf_vf_mux_scbd_174_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_174_up", this);
    pf_vf_mux_scbd_175_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_175_up", this);
    pf_vf_mux_scbd_176_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_176_up", this);
    pf_vf_mux_scbd_177_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_177_up", this);
    pf_vf_mux_scbd_178_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_178_up", this);
    pf_vf_mux_scbd_179_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_179_up", this);
    pf_vf_mux_scbd_180_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_180_up", this);
    pf_vf_mux_scbd_181_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_181_up", this);
    pf_vf_mux_scbd_182_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_182_up", this);
    pf_vf_mux_scbd_183_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_183_up", this);
    pf_vf_mux_scbd_184_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_184_up", this);
    pf_vf_mux_scbd_185_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_185_up", this);
    pf_vf_mux_scbd_186_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_186_up", this);
    pf_vf_mux_scbd_187_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_187_up", this);
    pf_vf_mux_scbd_188_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_188_up", this);
    pf_vf_mux_scbd_189_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_189_up", this);
    pf_vf_mux_scbd_190_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_190_up", this);
    pf_vf_mux_scbd_191_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_191_up", this);
    pf_vf_mux_scbd_192_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_192_up", this);
    pf_vf_mux_scbd_193_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_193_up", this);
    pf_vf_mux_scbd_194_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_194_up", this);
    pf_vf_mux_scbd_195_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_195_up", this);
    pf_vf_mux_scbd_196_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_196_up", this);
    pf_vf_mux_scbd_197_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_197_up", this);
    pf_vf_mux_scbd_198_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_198_up", this);
    pf_vf_mux_scbd_199_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_199_up", this);
    pf_vf_mux_scbd_200_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_200_up", this);
    pf_vf_mux_scbd_201_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_201_up", this);
    pf_vf_mux_scbd_202_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_202_up", this);
    pf_vf_mux_scbd_203_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_203_up", this);
    pf_vf_mux_scbd_204_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_204_up", this);
    pf_vf_mux_scbd_205_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_205_up", this);
    pf_vf_mux_scbd_206_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_206_up", this);
    pf_vf_mux_scbd_207_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_207_up", this);
    pf_vf_mux_scbd_208_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_208_up", this);
    pf_vf_mux_scbd_209_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_209_up", this);
    pf_vf_mux_scbd_210_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_210_up", this);
    pf_vf_mux_scbd_211_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_211_up", this);
    pf_vf_mux_scbd_212_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_212_up", this);
    pf_vf_mux_scbd_213_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_213_up", this);
    pf_vf_mux_scbd_214_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_214_up", this);
    pf_vf_mux_scbd_215_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_215_up", this);
    pf_vf_mux_scbd_216_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_216_up", this);
    pf_vf_mux_scbd_217_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_217_up", this);
    pf_vf_mux_scbd_218_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_218_up", this);
    pf_vf_mux_scbd_219_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_219_up", this);
    pf_vf_mux_scbd_220_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_220_up", this);
    pf_vf_mux_scbd_221_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_221_up", this);
    pf_vf_mux_scbd_222_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_222_up", this);
    pf_vf_mux_scbd_223_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_223_up", this);
    pf_vf_mux_scbd_224_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_224_up", this);
    pf_vf_mux_scbd_225_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_225_up", this);
    pf_vf_mux_scbd_226_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_226_up", this);
    pf_vf_mux_scbd_227_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_227_up", this);
    pf_vf_mux_scbd_228_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_228_up", this);
    pf_vf_mux_scbd_229_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_229_up", this);
    pf_vf_mux_scbd_230_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_230_up", this);
    pf_vf_mux_scbd_231_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_231_up", this);
    pf_vf_mux_scbd_232_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_232_up", this);
    pf_vf_mux_scbd_233_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_233_up", this);
    pf_vf_mux_scbd_234_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_234_up", this);
    pf_vf_mux_scbd_235_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_235_up", this);
    pf_vf_mux_scbd_236_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_236_up", this);
    pf_vf_mux_scbd_237_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_237_up", this);
    pf_vf_mux_scbd_238_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_238_up", this);
    pf_vf_mux_scbd_239_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_239_up", this);
    pf_vf_mux_scbd_240_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_240_up", this);
    pf_vf_mux_scbd_241_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_241_up", this);
    pf_vf_mux_scbd_242_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_242_up", this);
    pf_vf_mux_scbd_243_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_243_up", this);
    pf_vf_mux_scbd_244_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_244_up", this);
    pf_vf_mux_scbd_245_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_245_up", this);
    pf_vf_mux_scbd_246_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_246_up", this);
    pf_vf_mux_scbd_247_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_247_up", this);
    pf_vf_mux_scbd_248_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_248_up", this);
    pf_vf_mux_scbd_249_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_249_up", this);
    pf_vf_mux_scbd_250_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_250_up", this);
    pf_vf_mux_scbd_251_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_251_up", this);
    pf_vf_mux_scbd_252_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_252_up", this);
    pf_vf_mux_scbd_253_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_253_up", this);
    pf_vf_mux_scbd_254_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_254_up", this);
    pf_vf_mux_scbd_255_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_255_up", this);
    pf_vf_mux_scbd_256_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_256_up", this);
    pf_vf_mux_scbd_257_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_257_up", this);
    pf_vf_mux_scbd_258_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_258_up", this);
    pf_vf_mux_scbd_259_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_259_up", this);
    pf_vf_mux_scbd_260_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_260_up", this);
    pf_vf_mux_scbd_261_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_261_up", this);
    pf_vf_mux_scbd_262_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_262_up", this);
    pf_vf_mux_scbd_263_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_263_up", this);
    pf_vf_mux_scbd_264_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_264_up", this);
    pf_vf_mux_scbd_265_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_265_up", this);
    pf_vf_mux_scbd_266_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_266_up", this);
    pf_vf_mux_scbd_267_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_267_up", this);
    pf_vf_mux_scbd_268_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_268_up", this);
    pf_vf_mux_scbd_269_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_269_up", this);
    pf_vf_mux_scbd_270_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_270_up", this);
    pf_vf_mux_scbd_271_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_271_up", this);
    pf_vf_mux_scbd_272_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_272_up", this);
    pf_vf_mux_scbd_273_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_273_up", this);
    pf_vf_mux_scbd_274_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_274_up", this);
    pf_vf_mux_scbd_275_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_275_up", this);
    pf_vf_mux_scbd_276_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_276_up", this);
    pf_vf_mux_scbd_277_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_277_up", this);
    pf_vf_mux_scbd_278_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_278_up", this);
    pf_vf_mux_scbd_279_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_279_up", this);
    pf_vf_mux_scbd_280_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_280_up", this);
    pf_vf_mux_scbd_281_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_281_up", this);
    pf_vf_mux_scbd_282_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_282_up", this);
    pf_vf_mux_scbd_283_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_283_up", this);
    pf_vf_mux_scbd_284_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_284_up", this);
    pf_vf_mux_scbd_285_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_285_up", this);
    pf_vf_mux_scbd_286_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_286_up", this);
    pf_vf_mux_scbd_287_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_287_up", this);
    pf_vf_mux_scbd_288_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_288_up", this);
    pf_vf_mux_scbd_289_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_289_up", this);
    pf_vf_mux_scbd_290_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_290_up", this);
    pf_vf_mux_scbd_291_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_291_up", this);
    pf_vf_mux_scbd_292_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_292_up", this);
    pf_vf_mux_scbd_293_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_293_up", this);
    pf_vf_mux_scbd_294_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_294_up", this);
    pf_vf_mux_scbd_295_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_295_up", this);
    pf_vf_mux_scbd_296_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_296_up", this);
    pf_vf_mux_scbd_297_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_297_up", this);
    pf_vf_mux_scbd_298_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_298_up", this);
    pf_vf_mux_scbd_299_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_299_up", this);
    pf_vf_mux_scbd_300_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_300_up", this);
    pf_vf_mux_scbd_301_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_301_up", this);
    pf_vf_mux_scbd_302_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_302_up", this);
    pf_vf_mux_scbd_303_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_303_up", this);
    pf_vf_mux_scbd_304_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_304_up", this);
    pf_vf_mux_scbd_305_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_305_up", this);
    pf_vf_mux_scbd_306_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_306_up", this);
    pf_vf_mux_scbd_307_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_307_up", this);
    pf_vf_mux_scbd_308_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_308_up", this);
    pf_vf_mux_scbd_309_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_309_up", this);
    pf_vf_mux_scbd_310_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_310_up", this);
    pf_vf_mux_scbd_311_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_311_up", this);
    pf_vf_mux_scbd_312_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_312_up", this);
    pf_vf_mux_scbd_313_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_313_up", this);
    pf_vf_mux_scbd_314_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_314_up", this);
    pf_vf_mux_scbd_315_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_315_up", this);
    pf_vf_mux_scbd_316_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_316_up", this);
    pf_vf_mux_scbd_317_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_317_up", this);
    pf_vf_mux_scbd_318_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_318_up", this);
    pf_vf_mux_scbd_319_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_319_up", this);
    pf_vf_mux_scbd_320_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_320_up", this);
    pf_vf_mux_scbd_321_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_321_up", this);
    pf_vf_mux_scbd_322_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_322_up", this);
    pf_vf_mux_scbd_323_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_323_up", this);
    pf_vf_mux_scbd_324_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_324_up", this);
    pf_vf_mux_scbd_325_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_325_up", this);
    pf_vf_mux_scbd_326_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_326_up", this);
    pf_vf_mux_scbd_327_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_327_up", this);
    pf_vf_mux_scbd_328_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_328_up", this);
    pf_vf_mux_scbd_329_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_329_up", this);
    pf_vf_mux_scbd_330_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_330_up", this);
    pf_vf_mux_scbd_331_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_331_up", this);
    pf_vf_mux_scbd_332_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_332_up", this);
    pf_vf_mux_scbd_333_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_333_up", this);
    pf_vf_mux_scbd_334_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_334_up", this);
    pf_vf_mux_scbd_335_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_335_up", this);
    pf_vf_mux_scbd_336_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_336_up", this);
    pf_vf_mux_scbd_337_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_337_up", this);
    pf_vf_mux_scbd_338_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_338_up", this);
    pf_vf_mux_scbd_339_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_339_up", this);
    pf_vf_mux_scbd_340_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_340_up", this);
    pf_vf_mux_scbd_341_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_341_up", this);
    pf_vf_mux_scbd_342_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_342_up", this);
    pf_vf_mux_scbd_343_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_343_up", this);
    pf_vf_mux_scbd_344_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_344_up", this);
    pf_vf_mux_scbd_345_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_345_up", this);
    pf_vf_mux_scbd_346_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_346_up", this);
    pf_vf_mux_scbd_347_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_347_up", this);
    pf_vf_mux_scbd_348_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_348_up", this);
    pf_vf_mux_scbd_349_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_349_up", this);
    pf_vf_mux_scbd_350_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_350_up", this);
    pf_vf_mux_scbd_351_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_351_up", this);
    pf_vf_mux_scbd_352_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_352_up", this);
    pf_vf_mux_scbd_353_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_353_up", this);
    pf_vf_mux_scbd_354_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_354_up", this);
    pf_vf_mux_scbd_355_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_355_up", this);
    pf_vf_mux_scbd_356_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_356_up", this);
    pf_vf_mux_scbd_357_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_357_up", this);
    pf_vf_mux_scbd_358_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_358_up", this);
    pf_vf_mux_scbd_359_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_359_up", this);
    pf_vf_mux_scbd_360_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_360_up", this);
    pf_vf_mux_scbd_361_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_361_up", this);
    pf_vf_mux_scbd_362_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_362_up", this);
    pf_vf_mux_scbd_363_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_363_up", this);
    pf_vf_mux_scbd_364_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_364_up", this);
    pf_vf_mux_scbd_365_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_365_up", this);
    pf_vf_mux_scbd_366_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_366_up", this);
    pf_vf_mux_scbd_367_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_367_up", this);
    pf_vf_mux_scbd_368_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_368_up", this);
    pf_vf_mux_scbd_369_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_369_up", this);
    pf_vf_mux_scbd_370_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_370_up", this);
    pf_vf_mux_scbd_371_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_371_up", this);
    pf_vf_mux_scbd_372_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_372_up", this);
    pf_vf_mux_scbd_373_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_373_up", this);
    pf_vf_mux_scbd_374_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_374_up", this);
    pf_vf_mux_scbd_375_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_375_up", this);
    pf_vf_mux_scbd_376_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_376_up", this);
    pf_vf_mux_scbd_377_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_377_up", this);
    pf_vf_mux_scbd_378_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_378_up", this);
    pf_vf_mux_scbd_379_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_379_up", this);
    pf_vf_mux_scbd_380_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_380_up", this);
    pf_vf_mux_scbd_381_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_381_up", this);
    pf_vf_mux_scbd_382_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_382_up", this);
    pf_vf_mux_scbd_383_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_383_up", this);
    pf_vf_mux_scbd_384_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_384_up", this);
    pf_vf_mux_scbd_385_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_385_up", this);
    pf_vf_mux_scbd_386_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_386_up", this);
    pf_vf_mux_scbd_387_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_387_up", this);
    pf_vf_mux_scbd_388_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_388_up", this);
    pf_vf_mux_scbd_389_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_389_up", this);
    pf_vf_mux_scbd_390_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_390_up", this);
    pf_vf_mux_scbd_391_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_391_up", this);
    pf_vf_mux_scbd_392_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_392_up", this);
    pf_vf_mux_scbd_393_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_393_up", this);
    pf_vf_mux_scbd_394_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_394_up", this);
    pf_vf_mux_scbd_395_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_395_up", this);
    pf_vf_mux_scbd_396_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_396_up", this);
    pf_vf_mux_scbd_397_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_397_up", this);
    pf_vf_mux_scbd_398_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_398_up", this);
    pf_vf_mux_scbd_399_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_399_up", this);
    pf_vf_mux_scbd_400_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_400_up", this);
    pf_vf_mux_scbd_401_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_401_up", this);
    pf_vf_mux_scbd_402_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_402_up", this);
    pf_vf_mux_scbd_403_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_403_up", this);
    pf_vf_mux_scbd_404_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_404_up", this);
    pf_vf_mux_scbd_405_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_405_up", this);
    pf_vf_mux_scbd_406_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_406_up", this);
    pf_vf_mux_scbd_407_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_407_up", this);
    pf_vf_mux_scbd_408_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_408_up", this);
    pf_vf_mux_scbd_409_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_409_up", this);
    pf_vf_mux_scbd_410_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_410_up", this);
    pf_vf_mux_scbd_411_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_411_up", this);
    pf_vf_mux_scbd_412_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_412_up", this);
    pf_vf_mux_scbd_413_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_413_up", this);
    pf_vf_mux_scbd_414_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_414_up", this);
    pf_vf_mux_scbd_415_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_415_up", this);
    pf_vf_mux_scbd_416_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_416_up", this);
    pf_vf_mux_scbd_417_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_417_up", this);
    pf_vf_mux_scbd_418_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_418_up", this);
    pf_vf_mux_scbd_419_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_419_up", this);
    pf_vf_mux_scbd_420_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_420_up", this);
    pf_vf_mux_scbd_421_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_421_up", this);
    pf_vf_mux_scbd_422_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_422_up", this);
    pf_vf_mux_scbd_423_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_423_up", this);
    pf_vf_mux_scbd_424_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_424_up", this);
    pf_vf_mux_scbd_425_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_425_up", this);
    pf_vf_mux_scbd_426_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_426_up", this);
    pf_vf_mux_scbd_427_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_427_up", this);
    pf_vf_mux_scbd_428_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_428_up", this);
    pf_vf_mux_scbd_429_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_429_up", this);
    pf_vf_mux_scbd_430_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_430_up", this);
    pf_vf_mux_scbd_431_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_431_up", this);
    pf_vf_mux_scbd_432_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_432_up", this);
    pf_vf_mux_scbd_433_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_433_up", this);
    pf_vf_mux_scbd_434_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_434_up", this);
    pf_vf_mux_scbd_435_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_435_up", this);
    pf_vf_mux_scbd_436_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_436_up", this);
    pf_vf_mux_scbd_437_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_437_up", this);
    pf_vf_mux_scbd_438_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_438_up", this);
    pf_vf_mux_scbd_439_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_439_up", this);
    pf_vf_mux_scbd_440_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_440_up", this);
    pf_vf_mux_scbd_441_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_441_up", this);
    pf_vf_mux_scbd_442_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_442_up", this);
    pf_vf_mux_scbd_443_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_443_up", this);
    pf_vf_mux_scbd_444_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_444_up", this);
    pf_vf_mux_scbd_445_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_445_up", this);
    pf_vf_mux_scbd_446_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_446_up", this);
    pf_vf_mux_scbd_447_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_447_up", this);
    pf_vf_mux_scbd_448_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_448_up", this);
    pf_vf_mux_scbd_449_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_449_up", this);
    pf_vf_mux_scbd_450_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_450_up", this);
    pf_vf_mux_scbd_451_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_451_up", this);
    pf_vf_mux_scbd_452_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_452_up", this);
    pf_vf_mux_scbd_453_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_453_up", this);
    pf_vf_mux_scbd_454_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_454_up", this);
    pf_vf_mux_scbd_455_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_455_up", this);
    pf_vf_mux_scbd_456_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_456_up", this);
    pf_vf_mux_scbd_457_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_457_up", this);
    pf_vf_mux_scbd_458_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_458_up", this);
    pf_vf_mux_scbd_459_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_459_up", this);
    pf_vf_mux_scbd_460_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_460_up", this);
    pf_vf_mux_scbd_461_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_461_up", this);
    pf_vf_mux_scbd_462_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_462_up", this);
    pf_vf_mux_scbd_463_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_463_up", this);
    pf_vf_mux_scbd_464_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_464_up", this);
    pf_vf_mux_scbd_465_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_465_up", this);
    pf_vf_mux_scbd_466_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_466_up", this);
    pf_vf_mux_scbd_467_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_467_up", this);
    pf_vf_mux_scbd_468_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_468_up", this);
    pf_vf_mux_scbd_469_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_469_up", this);
    pf_vf_mux_scbd_470_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_470_up", this);
    pf_vf_mux_scbd_471_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_471_up", this);
    pf_vf_mux_scbd_472_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_472_up", this);
    pf_vf_mux_scbd_473_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_473_up", this);
    pf_vf_mux_scbd_474_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_474_up", this);
    pf_vf_mux_scbd_475_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_475_up", this);
    pf_vf_mux_scbd_476_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_476_up", this);
    pf_vf_mux_scbd_477_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_477_up", this);
    pf_vf_mux_scbd_478_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_478_up", this);
    pf_vf_mux_scbd_479_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_479_up", this);
    pf_vf_mux_scbd_480_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_480_up", this);
    pf_vf_mux_scbd_481_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_481_up", this);
    pf_vf_mux_scbd_482_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_482_up", this);
    pf_vf_mux_scbd_483_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_483_up", this);
    pf_vf_mux_scbd_484_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_484_up", this);
    pf_vf_mux_scbd_485_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_485_up", this);
    pf_vf_mux_scbd_486_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_486_up", this);
    pf_vf_mux_scbd_487_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_487_up", this);
    pf_vf_mux_scbd_488_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_488_up", this);
    pf_vf_mux_scbd_489_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_489_up", this);
    pf_vf_mux_scbd_490_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_490_up", this);
    pf_vf_mux_scbd_491_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_491_up", this);
    pf_vf_mux_scbd_492_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_492_up", this);
    pf_vf_mux_scbd_493_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_493_up", this);
    pf_vf_mux_scbd_494_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_494_up", this);
    pf_vf_mux_scbd_495_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_495_up", this);
    pf_vf_mux_scbd_496_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_496_up", this);
    pf_vf_mux_scbd_497_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_497_up", this);
    pf_vf_mux_scbd_498_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_498_up", this);
    pf_vf_mux_scbd_499_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_499_up", this);
    pf_vf_mux_scbd_500_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_500_up", this);
    pf_vf_mux_scbd_501_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_501_up", this);
    pf_vf_mux_scbd_502_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_502_up", this);
    pf_vf_mux_scbd_503_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_503_up", this);
    pf_vf_mux_scbd_504_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_504_up", this);
    pf_vf_mux_scbd_505_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_505_up", this);
    pf_vf_mux_scbd_506_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_506_up", this);
    pf_vf_mux_scbd_507_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_507_up", this);
    pf_vf_mux_scbd_508_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_508_up", this);
    pf_vf_mux_scbd_509_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_509_up", this);
    pf_vf_mux_scbd_510_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_510_up", this);
    pf_vf_mux_scbd_511_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_511_up", this);
    pf_vf_mux_scbd_512_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_512_up", this);
    pf_vf_mux_scbd_513_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_513_up", this);
    pf_vf_mux_scbd_514_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_514_up", this);
    pf_vf_mux_scbd_515_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_515_up", this);
    pf_vf_mux_scbd_516_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_516_up", this);
    pf_vf_mux_scbd_517_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_517_up", this);
    pf_vf_mux_scbd_518_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_518_up", this);
    pf_vf_mux_scbd_519_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_519_up", this);
    pf_vf_mux_scbd_520_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_520_up", this);
    pf_vf_mux_scbd_521_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_521_up", this);
    pf_vf_mux_scbd_522_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_522_up", this);
    pf_vf_mux_scbd_523_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_523_up", this);
    pf_vf_mux_scbd_524_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_524_up", this);
    pf_vf_mux_scbd_525_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_525_up", this);
    pf_vf_mux_scbd_526_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_526_up", this);
    pf_vf_mux_scbd_527_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_527_up", this);
    pf_vf_mux_scbd_528_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_528_up", this);
    pf_vf_mux_scbd_529_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_529_up", this);
    pf_vf_mux_scbd_530_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_530_up", this);
    pf_vf_mux_scbd_531_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_531_up", this);
    pf_vf_mux_scbd_532_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_532_up", this);
    pf_vf_mux_scbd_533_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_533_up", this);
    pf_vf_mux_scbd_534_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_534_up", this);
    pf_vf_mux_scbd_535_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_535_up", this);
    pf_vf_mux_scbd_536_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_536_up", this);
    pf_vf_mux_scbd_537_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_537_up", this);
    pf_vf_mux_scbd_538_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_538_up", this);
    pf_vf_mux_scbd_539_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_539_up", this);
    pf_vf_mux_scbd_540_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_540_up", this);
    pf_vf_mux_scbd_541_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_541_up", this);
    pf_vf_mux_scbd_542_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_542_up", this);
    pf_vf_mux_scbd_543_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_543_up", this);
    pf_vf_mux_scbd_544_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_544_up", this);
    pf_vf_mux_scbd_545_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_545_up", this);
    pf_vf_mux_scbd_546_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_546_up", this);
    pf_vf_mux_scbd_547_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_547_up", this);
    pf_vf_mux_scbd_548_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_548_up", this);
    pf_vf_mux_scbd_549_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_549_up", this);
    pf_vf_mux_scbd_550_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_550_up", this);
    pf_vf_mux_scbd_551_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_551_up", this);
    pf_vf_mux_scbd_552_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_552_up", this);
    pf_vf_mux_scbd_553_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_553_up", this);
    pf_vf_mux_scbd_554_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_554_up", this);
    pf_vf_mux_scbd_555_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_555_up", this);
    pf_vf_mux_scbd_556_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_556_up", this);
    pf_vf_mux_scbd_557_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_557_up", this);
    pf_vf_mux_scbd_558_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_558_up", this);
    pf_vf_mux_scbd_559_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_559_up", this);
    pf_vf_mux_scbd_560_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_560_up", this);
    pf_vf_mux_scbd_561_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_561_up", this);
    pf_vf_mux_scbd_562_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_562_up", this);
    pf_vf_mux_scbd_563_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_563_up", this);
    pf_vf_mux_scbd_564_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_564_up", this);
    pf_vf_mux_scbd_565_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_565_up", this);
    pf_vf_mux_scbd_566_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_566_up", this);
    pf_vf_mux_scbd_567_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_567_up", this);
    pf_vf_mux_scbd_568_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_568_up", this);
    pf_vf_mux_scbd_569_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_569_up", this);
    pf_vf_mux_scbd_570_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_570_up", this);
    pf_vf_mux_scbd_571_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_571_up", this);
    pf_vf_mux_scbd_572_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_572_up", this);
    pf_vf_mux_scbd_573_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_573_up", this);
    pf_vf_mux_scbd_574_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_574_up", this);
    pf_vf_mux_scbd_575_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_575_up", this);
    pf_vf_mux_scbd_576_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_576_up", this);
    pf_vf_mux_scbd_577_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_577_up", this);
    pf_vf_mux_scbd_578_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_578_up", this);
    pf_vf_mux_scbd_579_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_579_up", this);
    pf_vf_mux_scbd_580_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_580_up", this);
    pf_vf_mux_scbd_581_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_581_up", this);
    pf_vf_mux_scbd_582_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_582_up", this);
    pf_vf_mux_scbd_583_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_583_up", this);
    pf_vf_mux_scbd_584_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_584_up", this);
    pf_vf_mux_scbd_585_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_585_up", this);
    pf_vf_mux_scbd_586_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_586_up", this);
    pf_vf_mux_scbd_587_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_587_up", this);
    pf_vf_mux_scbd_588_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_588_up", this);
    pf_vf_mux_scbd_589_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_589_up", this);
    pf_vf_mux_scbd_590_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_590_up", this);
    pf_vf_mux_scbd_591_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_591_up", this);
    pf_vf_mux_scbd_592_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_592_up", this);
    pf_vf_mux_scbd_593_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_593_up", this);
    pf_vf_mux_scbd_594_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_594_up", this);
    pf_vf_mux_scbd_595_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_595_up", this);
    pf_vf_mux_scbd_596_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_596_up", this);
    pf_vf_mux_scbd_597_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_597_up", this);
    pf_vf_mux_scbd_598_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_598_up", this);
    pf_vf_mux_scbd_599_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_599_up", this);
    pf_vf_mux_scbd_600_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_600_up", this);
    pf_vf_mux_scbd_601_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_601_up", this);
    pf_vf_mux_scbd_602_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_602_up", this);
    pf_vf_mux_scbd_603_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_603_up", this);
    pf_vf_mux_scbd_604_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_604_up", this);
    pf_vf_mux_scbd_605_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_605_up", this);
    pf_vf_mux_scbd_606_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_606_up", this);
    pf_vf_mux_scbd_607_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_607_up", this);
    pf_vf_mux_scbd_608_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_608_up", this);
    pf_vf_mux_scbd_609_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_609_up", this);
    pf_vf_mux_scbd_610_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_610_up", this);
    pf_vf_mux_scbd_611_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_611_up", this);
    pf_vf_mux_scbd_612_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_612_up", this);
    pf_vf_mux_scbd_613_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_613_up", this);
    pf_vf_mux_scbd_614_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_614_up", this);
    pf_vf_mux_scbd_615_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_615_up", this);
    pf_vf_mux_scbd_616_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_616_up", this);
    pf_vf_mux_scbd_617_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_617_up", this);
    pf_vf_mux_scbd_618_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_618_up", this);
    pf_vf_mux_scbd_619_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_619_up", this);
    pf_vf_mux_scbd_620_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_620_up", this);
    pf_vf_mux_scbd_621_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_621_up", this);
    pf_vf_mux_scbd_622_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_622_up", this);
    pf_vf_mux_scbd_623_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_623_up", this);
    pf_vf_mux_scbd_624_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_624_up", this);
    pf_vf_mux_scbd_625_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_625_up", this);
    pf_vf_mux_scbd_626_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_626_up", this);
    pf_vf_mux_scbd_627_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_627_up", this);
    pf_vf_mux_scbd_628_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_628_up", this);
    pf_vf_mux_scbd_629_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_629_up", this);
    pf_vf_mux_scbd_630_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_630_up", this);
    pf_vf_mux_scbd_631_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_631_up", this);
    pf_vf_mux_scbd_632_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_632_up", this);
    pf_vf_mux_scbd_633_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_633_up", this);
    pf_vf_mux_scbd_634_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_634_up", this);
    pf_vf_mux_scbd_635_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_635_up", this);
    pf_vf_mux_scbd_636_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_636_up", this);
    pf_vf_mux_scbd_637_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_637_up", this);
    pf_vf_mux_scbd_638_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_638_up", this);
    pf_vf_mux_scbd_639_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_639_up", this);
    pf_vf_mux_scbd_640_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_640_up", this);
    pf_vf_mux_scbd_641_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_641_up", this);
    pf_vf_mux_scbd_642_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_642_up", this);
    pf_vf_mux_scbd_643_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_643_up", this);
    pf_vf_mux_scbd_644_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_644_up", this);
    pf_vf_mux_scbd_645_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_645_up", this);
    pf_vf_mux_scbd_646_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_646_up", this);
    pf_vf_mux_scbd_647_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_647_up", this);
    pf_vf_mux_scbd_648_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_648_up", this);
    pf_vf_mux_scbd_649_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_649_up", this);
    pf_vf_mux_scbd_650_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_650_up", this);
    pf_vf_mux_scbd_651_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_651_up", this);
    pf_vf_mux_scbd_652_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_652_up", this);
    pf_vf_mux_scbd_653_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_653_up", this);
    pf_vf_mux_scbd_654_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_654_up", this);
    pf_vf_mux_scbd_655_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_655_up", this);
    pf_vf_mux_scbd_656_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_656_up", this);
    pf_vf_mux_scbd_657_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_657_up", this);
    pf_vf_mux_scbd_658_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_658_up", this);
    pf_vf_mux_scbd_659_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_659_up", this);
    pf_vf_mux_scbd_660_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_660_up", this);
    pf_vf_mux_scbd_661_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_661_up", this);
    pf_vf_mux_scbd_662_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_662_up", this);
    pf_vf_mux_scbd_663_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_663_up", this);
    pf_vf_mux_scbd_664_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_664_up", this);
    pf_vf_mux_scbd_665_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_665_up", this);
    pf_vf_mux_scbd_666_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_666_up", this);
    pf_vf_mux_scbd_667_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_667_up", this);
    pf_vf_mux_scbd_668_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_668_up", this);
    pf_vf_mux_scbd_669_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_669_up", this);
    pf_vf_mux_scbd_670_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_670_up", this);
    pf_vf_mux_scbd_671_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_671_up", this);
    pf_vf_mux_scbd_672_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_672_up", this);
    pf_vf_mux_scbd_673_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_673_up", this);
    pf_vf_mux_scbd_674_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_674_up", this);
    pf_vf_mux_scbd_675_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_675_up", this);
    pf_vf_mux_scbd_676_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_676_up", this);
    pf_vf_mux_scbd_677_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_677_up", this);
    pf_vf_mux_scbd_678_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_678_up", this);
    pf_vf_mux_scbd_679_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_679_up", this);
    pf_vf_mux_scbd_680_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_680_up", this);
    pf_vf_mux_scbd_681_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_681_up", this);
    pf_vf_mux_scbd_682_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_682_up", this);
    pf_vf_mux_scbd_683_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_683_up", this);
    pf_vf_mux_scbd_684_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_684_up", this);
    pf_vf_mux_scbd_685_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_685_up", this);
    pf_vf_mux_scbd_686_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_686_up", this);
    pf_vf_mux_scbd_687_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_687_up", this);
    pf_vf_mux_scbd_688_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_688_up", this);
    pf_vf_mux_scbd_689_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_689_up", this);
    pf_vf_mux_scbd_690_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_690_up", this);
    pf_vf_mux_scbd_691_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_691_up", this);
    pf_vf_mux_scbd_692_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_692_up", this);
    pf_vf_mux_scbd_693_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_693_up", this);
    pf_vf_mux_scbd_694_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_694_up", this);
    pf_vf_mux_scbd_695_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_695_up", this);
    pf_vf_mux_scbd_696_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_696_up", this);
    pf_vf_mux_scbd_697_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_697_up", this);
    pf_vf_mux_scbd_698_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_698_up", this);
    pf_vf_mux_scbd_699_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_699_up", this);
    pf_vf_mux_scbd_700_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_700_up", this);
    pf_vf_mux_scbd_701_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_701_up", this);
    pf_vf_mux_scbd_702_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_702_up", this);
    pf_vf_mux_scbd_703_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_703_up", this);
    pf_vf_mux_scbd_704_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_704_up", this);
    pf_vf_mux_scbd_705_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_705_up", this);
    pf_vf_mux_scbd_706_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_706_up", this);
    pf_vf_mux_scbd_707_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_707_up", this);
    pf_vf_mux_scbd_708_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_708_up", this);
    pf_vf_mux_scbd_709_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_709_up", this);
    pf_vf_mux_scbd_710_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_710_up", this);
    pf_vf_mux_scbd_711_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_711_up", this);
    pf_vf_mux_scbd_712_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_712_up", this);
    pf_vf_mux_scbd_713_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_713_up", this);
    pf_vf_mux_scbd_714_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_714_up", this);
    pf_vf_mux_scbd_715_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_715_up", this);
    pf_vf_mux_scbd_716_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_716_up", this);
    pf_vf_mux_scbd_717_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_717_up", this);
    pf_vf_mux_scbd_718_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_718_up", this);
    pf_vf_mux_scbd_719_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_719_up", this);
    pf_vf_mux_scbd_720_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_720_up", this);
    pf_vf_mux_scbd_721_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_721_up", this);
    pf_vf_mux_scbd_722_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_722_up", this);
    pf_vf_mux_scbd_723_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_723_up", this);
    pf_vf_mux_scbd_724_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_724_up", this);
    pf_vf_mux_scbd_725_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_725_up", this);
    pf_vf_mux_scbd_726_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_726_up", this);
    pf_vf_mux_scbd_727_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_727_up", this);
    pf_vf_mux_scbd_728_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_728_up", this);
    pf_vf_mux_scbd_729_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_729_up", this);
    pf_vf_mux_scbd_730_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_730_up", this);
    pf_vf_mux_scbd_731_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_731_up", this);
    pf_vf_mux_scbd_732_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_732_up", this);
    pf_vf_mux_scbd_733_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_733_up", this);
    pf_vf_mux_scbd_734_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_734_up", this);
    pf_vf_mux_scbd_735_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_735_up", this);
    pf_vf_mux_scbd_736_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_736_up", this);
    pf_vf_mux_scbd_737_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_737_up", this);
    pf_vf_mux_scbd_738_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_738_up", this);
    pf_vf_mux_scbd_739_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_739_up", this);
    pf_vf_mux_scbd_740_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_740_up", this);
    pf_vf_mux_scbd_741_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_741_up", this);
    pf_vf_mux_scbd_742_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_742_up", this);
    pf_vf_mux_scbd_743_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_743_up", this);
    pf_vf_mux_scbd_744_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_744_up", this);
    pf_vf_mux_scbd_745_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_745_up", this);
    pf_vf_mux_scbd_746_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_746_up", this);
    pf_vf_mux_scbd_747_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_747_up", this);
    pf_vf_mux_scbd_748_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_748_up", this);
    pf_vf_mux_scbd_749_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_749_up", this);
    pf_vf_mux_scbd_750_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_750_up", this);
    pf_vf_mux_scbd_751_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_751_up", this);
    pf_vf_mux_scbd_752_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_752_up", this);
    pf_vf_mux_scbd_753_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_753_up", this);
    pf_vf_mux_scbd_754_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_754_up", this);
    pf_vf_mux_scbd_755_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_755_up", this);
    pf_vf_mux_scbd_756_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_756_up", this);
    pf_vf_mux_scbd_757_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_757_up", this);
    pf_vf_mux_scbd_758_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_758_up", this);
    pf_vf_mux_scbd_759_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_759_up", this);
    pf_vf_mux_scbd_760_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_760_up", this);
    pf_vf_mux_scbd_761_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_761_up", this);
    pf_vf_mux_scbd_762_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_762_up", this);
    pf_vf_mux_scbd_763_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_763_up", this);
    pf_vf_mux_scbd_764_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_764_up", this);
    pf_vf_mux_scbd_765_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_765_up", this);
    pf_vf_mux_scbd_766_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_766_up", this);
    pf_vf_mux_scbd_767_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_767_up", this);
    pf_vf_mux_scbd_768_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_768_up", this);
    pf_vf_mux_scbd_769_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_769_up", this);
    pf_vf_mux_scbd_770_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_770_up", this);
    pf_vf_mux_scbd_771_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_771_up", this);
    pf_vf_mux_scbd_772_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_772_up", this);
    pf_vf_mux_scbd_773_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_773_up", this);
    pf_vf_mux_scbd_774_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_774_up", this);
    pf_vf_mux_scbd_775_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_775_up", this);
    pf_vf_mux_scbd_776_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_776_up", this);
    pf_vf_mux_scbd_777_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_777_up", this);
    pf_vf_mux_scbd_778_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_778_up", this);
    pf_vf_mux_scbd_779_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_779_up", this);
    pf_vf_mux_scbd_780_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_780_up", this);
    pf_vf_mux_scbd_781_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_781_up", this);
    pf_vf_mux_scbd_782_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_782_up", this);
    pf_vf_mux_scbd_783_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_783_up", this);
    pf_vf_mux_scbd_784_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_784_up", this);
    pf_vf_mux_scbd_785_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_785_up", this);
    pf_vf_mux_scbd_786_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_786_up", this);
    pf_vf_mux_scbd_787_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_787_up", this);
    pf_vf_mux_scbd_788_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_788_up", this);
    pf_vf_mux_scbd_789_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_789_up", this);
    pf_vf_mux_scbd_790_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_790_up", this);
    pf_vf_mux_scbd_791_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_791_up", this);
    pf_vf_mux_scbd_792_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_792_up", this);
    pf_vf_mux_scbd_793_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_793_up", this);
    pf_vf_mux_scbd_794_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_794_up", this);
    pf_vf_mux_scbd_795_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_795_up", this);
    pf_vf_mux_scbd_796_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_796_up", this);
    pf_vf_mux_scbd_797_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_797_up", this);
    pf_vf_mux_scbd_798_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_798_up", this);
    pf_vf_mux_scbd_799_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_799_up", this);
    pf_vf_mux_scbd_800_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_800_up", this);
    pf_vf_mux_scbd_801_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_801_up", this);
    pf_vf_mux_scbd_802_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_802_up", this);
    pf_vf_mux_scbd_803_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_803_up", this);
    pf_vf_mux_scbd_804_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_804_up", this);
    pf_vf_mux_scbd_805_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_805_up", this);
    pf_vf_mux_scbd_806_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_806_up", this);
    pf_vf_mux_scbd_807_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_807_up", this);
    pf_vf_mux_scbd_808_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_808_up", this);
    pf_vf_mux_scbd_809_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_809_up", this);
    pf_vf_mux_scbd_810_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_810_up", this);
    pf_vf_mux_scbd_811_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_811_up", this);
    pf_vf_mux_scbd_812_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_812_up", this);
    pf_vf_mux_scbd_813_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_813_up", this);
    pf_vf_mux_scbd_814_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_814_up", this);
    pf_vf_mux_scbd_815_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_815_up", this);
    pf_vf_mux_scbd_816_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_816_up", this);
    pf_vf_mux_scbd_817_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_817_up", this);
    pf_vf_mux_scbd_818_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_818_up", this);
    pf_vf_mux_scbd_819_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_819_up", this);
    pf_vf_mux_scbd_820_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_820_up", this);
    pf_vf_mux_scbd_821_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_821_up", this);
    pf_vf_mux_scbd_822_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_822_up", this);
    pf_vf_mux_scbd_823_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_823_up", this);
    pf_vf_mux_scbd_824_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_824_up", this);
    pf_vf_mux_scbd_825_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_825_up", this);
    pf_vf_mux_scbd_826_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_826_up", this);
    pf_vf_mux_scbd_827_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_827_up", this);
    pf_vf_mux_scbd_828_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_828_up", this);
    pf_vf_mux_scbd_829_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_829_up", this);
    pf_vf_mux_scbd_830_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_830_up", this);
    pf_vf_mux_scbd_831_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_831_up", this);
    pf_vf_mux_scbd_832_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_832_up", this);
    pf_vf_mux_scbd_833_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_833_up", this);
    pf_vf_mux_scbd_834_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_834_up", this);
    pf_vf_mux_scbd_835_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_835_up", this);
    pf_vf_mux_scbd_836_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_836_up", this);
    pf_vf_mux_scbd_837_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_837_up", this);
    pf_vf_mux_scbd_838_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_838_up", this);
    pf_vf_mux_scbd_839_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_839_up", this);
    pf_vf_mux_scbd_840_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_840_up", this);
    pf_vf_mux_scbd_841_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_841_up", this);
    pf_vf_mux_scbd_842_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_842_up", this);
    pf_vf_mux_scbd_843_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_843_up", this);
    pf_vf_mux_scbd_844_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_844_up", this);
    pf_vf_mux_scbd_845_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_845_up", this);
    pf_vf_mux_scbd_846_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_846_up", this);
    pf_vf_mux_scbd_847_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_847_up", this);
    pf_vf_mux_scbd_848_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_848_up", this);
    pf_vf_mux_scbd_849_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_849_up", this);
    pf_vf_mux_scbd_850_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_850_up", this);
    pf_vf_mux_scbd_851_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_851_up", this);
    pf_vf_mux_scbd_852_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_852_up", this);
    pf_vf_mux_scbd_853_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_853_up", this);
    pf_vf_mux_scbd_854_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_854_up", this);
    pf_vf_mux_scbd_855_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_855_up", this);
    pf_vf_mux_scbd_856_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_856_up", this);
    pf_vf_mux_scbd_857_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_857_up", this);
    pf_vf_mux_scbd_858_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_858_up", this);
    pf_vf_mux_scbd_859_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_859_up", this);
    pf_vf_mux_scbd_860_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_860_up", this);
    pf_vf_mux_scbd_861_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_861_up", this);
    pf_vf_mux_scbd_862_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_862_up", this);
    pf_vf_mux_scbd_863_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_863_up", this);
    pf_vf_mux_scbd_864_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_864_up", this);
    pf_vf_mux_scbd_865_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_865_up", this);
    pf_vf_mux_scbd_866_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_866_up", this);
    pf_vf_mux_scbd_867_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_867_up", this);
    pf_vf_mux_scbd_868_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_868_up", this);
    pf_vf_mux_scbd_869_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_869_up", this);
    pf_vf_mux_scbd_870_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_870_up", this);
    pf_vf_mux_scbd_871_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_871_up", this);
    pf_vf_mux_scbd_872_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_872_up", this);
    pf_vf_mux_scbd_873_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_873_up", this);
    pf_vf_mux_scbd_874_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_874_up", this);
    pf_vf_mux_scbd_875_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_875_up", this);
    pf_vf_mux_scbd_876_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_876_up", this);
    pf_vf_mux_scbd_877_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_877_up", this);
    pf_vf_mux_scbd_878_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_878_up", this);
    pf_vf_mux_scbd_879_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_879_up", this);
    pf_vf_mux_scbd_880_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_880_up", this);
    pf_vf_mux_scbd_881_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_881_up", this);
    pf_vf_mux_scbd_882_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_882_up", this);
    pf_vf_mux_scbd_883_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_883_up", this);
    pf_vf_mux_scbd_884_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_884_up", this);
    pf_vf_mux_scbd_885_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_885_up", this);
    pf_vf_mux_scbd_886_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_886_up", this);
    pf_vf_mux_scbd_887_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_887_up", this);
    pf_vf_mux_scbd_888_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_888_up", this);
    pf_vf_mux_scbd_889_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_889_up", this);
    pf_vf_mux_scbd_890_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_890_up", this);
    pf_vf_mux_scbd_891_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_891_up", this);
    pf_vf_mux_scbd_892_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_892_up", this);
    pf_vf_mux_scbd_893_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_893_up", this);
    pf_vf_mux_scbd_894_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_894_up", this);
    pf_vf_mux_scbd_895_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_895_up", this);
    pf_vf_mux_scbd_896_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_896_up", this);
    pf_vf_mux_scbd_897_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_897_up", this);
    pf_vf_mux_scbd_898_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_898_up", this);
    pf_vf_mux_scbd_899_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_899_up", this);
    pf_vf_mux_scbd_900_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_900_up", this);
    pf_vf_mux_scbd_901_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_901_up", this);
    pf_vf_mux_scbd_902_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_902_up", this);
    pf_vf_mux_scbd_903_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_903_up", this);
    pf_vf_mux_scbd_904_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_904_up", this);
    pf_vf_mux_scbd_905_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_905_up", this);
    pf_vf_mux_scbd_906_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_906_up", this);
    pf_vf_mux_scbd_907_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_907_up", this);
    pf_vf_mux_scbd_908_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_908_up", this);
    pf_vf_mux_scbd_909_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_909_up", this);
    pf_vf_mux_scbd_910_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_910_up", this);
    pf_vf_mux_scbd_911_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_911_up", this);
    pf_vf_mux_scbd_912_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_912_up", this);
    pf_vf_mux_scbd_913_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_913_up", this);
    pf_vf_mux_scbd_914_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_914_up", this);
    pf_vf_mux_scbd_915_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_915_up", this);
    pf_vf_mux_scbd_916_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_916_up", this);
    pf_vf_mux_scbd_917_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_917_up", this);
    pf_vf_mux_scbd_918_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_918_up", this);
    pf_vf_mux_scbd_919_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_919_up", this);
    pf_vf_mux_scbd_920_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_920_up", this);
    pf_vf_mux_scbd_921_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_921_up", this);
    pf_vf_mux_scbd_922_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_922_up", this);
    pf_vf_mux_scbd_923_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_923_up", this);
    pf_vf_mux_scbd_924_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_924_up", this);
    pf_vf_mux_scbd_925_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_925_up", this);
    pf_vf_mux_scbd_926_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_926_up", this);
    pf_vf_mux_scbd_927_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_927_up", this);
    pf_vf_mux_scbd_928_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_928_up", this);
    pf_vf_mux_scbd_929_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_929_up", this);
    pf_vf_mux_scbd_930_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_930_up", this);
    pf_vf_mux_scbd_931_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_931_up", this);
    pf_vf_mux_scbd_932_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_932_up", this);
    pf_vf_mux_scbd_933_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_933_up", this);
    pf_vf_mux_scbd_934_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_934_up", this);
    pf_vf_mux_scbd_935_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_935_up", this);
    pf_vf_mux_scbd_936_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_936_up", this);
    pf_vf_mux_scbd_937_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_937_up", this);
    pf_vf_mux_scbd_938_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_938_up", this);
    pf_vf_mux_scbd_939_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_939_up", this);
    pf_vf_mux_scbd_940_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_940_up", this);
    pf_vf_mux_scbd_941_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_941_up", this);
    pf_vf_mux_scbd_942_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_942_up", this);
    pf_vf_mux_scbd_943_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_943_up", this);
    pf_vf_mux_scbd_944_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_944_up", this);
    pf_vf_mux_scbd_945_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_945_up", this);
    pf_vf_mux_scbd_946_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_946_up", this);
    pf_vf_mux_scbd_947_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_947_up", this);
    pf_vf_mux_scbd_948_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_948_up", this);
    pf_vf_mux_scbd_949_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_949_up", this);
    pf_vf_mux_scbd_950_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_950_up", this);
    pf_vf_mux_scbd_951_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_951_up", this);
    pf_vf_mux_scbd_952_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_952_up", this);
    pf_vf_mux_scbd_953_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_953_up", this);
    pf_vf_mux_scbd_954_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_954_up", this);
    pf_vf_mux_scbd_955_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_955_up", this);
    pf_vf_mux_scbd_956_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_956_up", this);
    pf_vf_mux_scbd_957_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_957_up", this);
    pf_vf_mux_scbd_958_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_958_up", this);
    pf_vf_mux_scbd_959_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_959_up", this);
    pf_vf_mux_scbd_960_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_960_up", this);
    pf_vf_mux_scbd_961_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_961_up", this);
    pf_vf_mux_scbd_962_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_962_up", this);
    pf_vf_mux_scbd_963_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_963_up", this);
    pf_vf_mux_scbd_964_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_964_up", this);
    pf_vf_mux_scbd_965_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_965_up", this);
    pf_vf_mux_scbd_966_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_966_up", this);
    pf_vf_mux_scbd_967_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_967_up", this);
    pf_vf_mux_scbd_968_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_968_up", this);
    pf_vf_mux_scbd_969_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_969_up", this);
    pf_vf_mux_scbd_970_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_970_up", this);
    pf_vf_mux_scbd_971_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_971_up", this);
    pf_vf_mux_scbd_972_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_972_up", this);
    pf_vf_mux_scbd_973_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_973_up", this);
    pf_vf_mux_scbd_974_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_974_up", this);
    pf_vf_mux_scbd_975_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_975_up", this);
    pf_vf_mux_scbd_976_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_976_up", this);
    pf_vf_mux_scbd_977_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_977_up", this);
    pf_vf_mux_scbd_978_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_978_up", this);
    pf_vf_mux_scbd_979_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_979_up", this);
    pf_vf_mux_scbd_980_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_980_up", this);
    pf_vf_mux_scbd_981_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_981_up", this);
    pf_vf_mux_scbd_982_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_982_up", this);
    pf_vf_mux_scbd_983_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_983_up", this);
    pf_vf_mux_scbd_984_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_984_up", this);
    pf_vf_mux_scbd_985_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_985_up", this);
    pf_vf_mux_scbd_986_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_986_up", this);
    pf_vf_mux_scbd_987_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_987_up", this);
    pf_vf_mux_scbd_988_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_988_up", this);
    pf_vf_mux_scbd_989_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_989_up", this);
    pf_vf_mux_scbd_990_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_990_up", this);
    pf_vf_mux_scbd_991_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_991_up", this);
    pf_vf_mux_scbd_992_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_992_up", this);
    pf_vf_mux_scbd_993_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_993_up", this);
    pf_vf_mux_scbd_994_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_994_up", this);
    pf_vf_mux_scbd_995_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_995_up", this);
    pf_vf_mux_scbd_996_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_996_up", this);
    pf_vf_mux_scbd_997_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_997_up", this);
    pf_vf_mux_scbd_998_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_998_up", this);
    pf_vf_mux_scbd_999_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_999_up", this);
    pf_vf_mux_scbd_1000_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1000_up", this);
    pf_vf_mux_scbd_1001_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1001_up", this);
    pf_vf_mux_scbd_1002_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1002_up", this);
    pf_vf_mux_scbd_1003_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1003_up", this);
    pf_vf_mux_scbd_1004_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1004_up", this);
    pf_vf_mux_scbd_1005_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1005_up", this);
    pf_vf_mux_scbd_1006_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1006_up", this);
    pf_vf_mux_scbd_1007_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1007_up", this);
    pf_vf_mux_scbd_1008_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1008_up", this);
    pf_vf_mux_scbd_1009_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1009_up", this);
    pf_vf_mux_scbd_1010_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1010_up", this);
    pf_vf_mux_scbd_1011_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1011_up", this);
    pf_vf_mux_scbd_1012_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1012_up", this);
    pf_vf_mux_scbd_1013_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1013_up", this);
    pf_vf_mux_scbd_1014_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1014_up", this);
    pf_vf_mux_scbd_1015_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1015_up", this);
    pf_vf_mux_scbd_1016_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1016_up", this);
    pf_vf_mux_scbd_1017_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1017_up", this);
    pf_vf_mux_scbd_1018_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1018_up", this);
    pf_vf_mux_scbd_1019_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1019_up", this);
    pf_vf_mux_scbd_1020_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1020_up", this);
    pf_vf_mux_scbd_1021_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1021_up", this);
    pf_vf_mux_scbd_1022_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1022_up", this);
    pf_vf_mux_scbd_1023_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1023_up", this);
    pf_vf_mux_scbd_1024_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1024_up", this);
    pf_vf_mux_scbd_1025_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1025_up", this);
    pf_vf_mux_scbd_1026_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1026_up", this);
    pf_vf_mux_scbd_1027_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1027_up", this);
    pf_vf_mux_scbd_1028_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1028_up", this);
    pf_vf_mux_scbd_1029_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1029_up", this);
    pf_vf_mux_scbd_1030_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1030_up", this);
    pf_vf_mux_scbd_1031_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1031_up", this);
    pf_vf_mux_scbd_1032_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1032_up", this);
    pf_vf_mux_scbd_1033_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1033_up", this);
    pf_vf_mux_scbd_1034_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1034_up", this);
    pf_vf_mux_scbd_1035_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1035_up", this);
    pf_vf_mux_scbd_1036_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1036_up", this);
    pf_vf_mux_scbd_1037_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1037_up", this);
    pf_vf_mux_scbd_1038_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1038_up", this);
    pf_vf_mux_scbd_1039_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1039_up", this);
    pf_vf_mux_scbd_1040_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1040_up", this);
    pf_vf_mux_scbd_1041_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1041_up", this);
    pf_vf_mux_scbd_1042_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1042_up", this);
    pf_vf_mux_scbd_1043_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1043_up", this);
    pf_vf_mux_scbd_1044_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1044_up", this);
    pf_vf_mux_scbd_1045_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1045_up", this);
    pf_vf_mux_scbd_1046_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1046_up", this);
    pf_vf_mux_scbd_1047_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1047_up", this);
    pf_vf_mux_scbd_1048_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1048_up", this);
    pf_vf_mux_scbd_1049_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1049_up", this);
    pf_vf_mux_scbd_1050_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1050_up", this);
    pf_vf_mux_scbd_1051_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1051_up", this);
    pf_vf_mux_scbd_1052_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1052_up", this);
    pf_vf_mux_scbd_1053_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1053_up", this);
    pf_vf_mux_scbd_1054_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1054_up", this);
    pf_vf_mux_scbd_1055_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1055_up", this);
    pf_vf_mux_scbd_1056_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1056_up", this);
    pf_vf_mux_scbd_1057_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1057_up", this);
    pf_vf_mux_scbd_1058_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1058_up", this);
    pf_vf_mux_scbd_1059_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1059_up", this);
    pf_vf_mux_scbd_1060_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1060_up", this);
    pf_vf_mux_scbd_1061_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1061_up", this);
    pf_vf_mux_scbd_1062_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1062_up", this);
    pf_vf_mux_scbd_1063_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1063_up", this);
    pf_vf_mux_scbd_1064_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1064_up", this);
    pf_vf_mux_scbd_1065_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1065_up", this);
    pf_vf_mux_scbd_1066_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1066_up", this);
    pf_vf_mux_scbd_1067_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1067_up", this);
    pf_vf_mux_scbd_1068_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1068_up", this);
    pf_vf_mux_scbd_1069_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1069_up", this);
    pf_vf_mux_scbd_1070_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1070_up", this);
    pf_vf_mux_scbd_1071_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1071_up", this);
    pf_vf_mux_scbd_1072_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1072_up", this);
    pf_vf_mux_scbd_1073_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1073_up", this);
    pf_vf_mux_scbd_1074_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1074_up", this);
    pf_vf_mux_scbd_1075_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1075_up", this);
    pf_vf_mux_scbd_1076_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1076_up", this);
    pf_vf_mux_scbd_1077_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1077_up", this);
    pf_vf_mux_scbd_1078_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1078_up", this);
    pf_vf_mux_scbd_1079_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1079_up", this);
    pf_vf_mux_scbd_1080_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1080_up", this);
    pf_vf_mux_scbd_1081_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1081_up", this);
    pf_vf_mux_scbd_1082_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1082_up", this);
    pf_vf_mux_scbd_1083_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1083_up", this);
    pf_vf_mux_scbd_1084_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1084_up", this);
    pf_vf_mux_scbd_1085_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1085_up", this);
    pf_vf_mux_scbd_1086_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1086_up", this);
    pf_vf_mux_scbd_1087_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1087_up", this);
    pf_vf_mux_scbd_1088_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1088_up", this);
    pf_vf_mux_scbd_1089_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1089_up", this);
    pf_vf_mux_scbd_1090_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1090_up", this);
    pf_vf_mux_scbd_1091_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1091_up", this);
    pf_vf_mux_scbd_1092_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1092_up", this);
    pf_vf_mux_scbd_1093_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1093_up", this);
    pf_vf_mux_scbd_1094_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1094_up", this);
    pf_vf_mux_scbd_1095_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1095_up", this);
    pf_vf_mux_scbd_1096_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1096_up", this);
    pf_vf_mux_scbd_1097_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1097_up", this);
    pf_vf_mux_scbd_1098_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1098_up", this);
    pf_vf_mux_scbd_1099_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1099_up", this);
    pf_vf_mux_scbd_1100_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1100_up", this);
    pf_vf_mux_scbd_1101_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1101_up", this);
    pf_vf_mux_scbd_1102_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1102_up", this);
    pf_vf_mux_scbd_1103_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1103_up", this);
    pf_vf_mux_scbd_1104_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1104_up", this);
    pf_vf_mux_scbd_1105_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1105_up", this);
    pf_vf_mux_scbd_1106_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1106_up", this);
    pf_vf_mux_scbd_1107_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1107_up", this);
    pf_vf_mux_scbd_1108_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1108_up", this);
    pf_vf_mux_scbd_1109_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1109_up", this);
    pf_vf_mux_scbd_1110_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1110_up", this);
    pf_vf_mux_scbd_1111_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1111_up", this);
    pf_vf_mux_scbd_1112_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1112_up", this);
    pf_vf_mux_scbd_1113_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1113_up", this);
    pf_vf_mux_scbd_1114_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1114_up", this);
    pf_vf_mux_scbd_1115_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1115_up", this);
    pf_vf_mux_scbd_1116_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1116_up", this);
    pf_vf_mux_scbd_1117_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1117_up", this);
    pf_vf_mux_scbd_1118_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1118_up", this);
    pf_vf_mux_scbd_1119_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1119_up", this);
    pf_vf_mux_scbd_1120_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1120_up", this);
    pf_vf_mux_scbd_1121_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1121_up", this);
    pf_vf_mux_scbd_1122_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1122_up", this);
    pf_vf_mux_scbd_1123_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1123_up", this);
    pf_vf_mux_scbd_1124_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1124_up", this);
    pf_vf_mux_scbd_1125_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1125_up", this);
    pf_vf_mux_scbd_1126_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1126_up", this);
    pf_vf_mux_scbd_1127_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1127_up", this);
    pf_vf_mux_scbd_1128_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1128_up", this);
    pf_vf_mux_scbd_1129_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1129_up", this);
    pf_vf_mux_scbd_1130_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1130_up", this);
    pf_vf_mux_scbd_1131_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1131_up", this);
    pf_vf_mux_scbd_1132_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1132_up", this);
    pf_vf_mux_scbd_1133_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1133_up", this);
    pf_vf_mux_scbd_1134_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1134_up", this);
    pf_vf_mux_scbd_1135_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1135_up", this);
    pf_vf_mux_scbd_1136_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1136_up", this);
    pf_vf_mux_scbd_1137_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1137_up", this);
    pf_vf_mux_scbd_1138_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1138_up", this);
    pf_vf_mux_scbd_1139_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1139_up", this);
    pf_vf_mux_scbd_1140_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1140_up", this);
    pf_vf_mux_scbd_1141_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1141_up", this);
    pf_vf_mux_scbd_1142_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1142_up", this);
    pf_vf_mux_scbd_1143_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1143_up", this);
    pf_vf_mux_scbd_1144_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1144_up", this);
    pf_vf_mux_scbd_1145_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1145_up", this);
    pf_vf_mux_scbd_1146_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1146_up", this);
    pf_vf_mux_scbd_1147_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1147_up", this);
    pf_vf_mux_scbd_1148_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1148_up", this);
    pf_vf_mux_scbd_1149_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1149_up", this);
    pf_vf_mux_scbd_1150_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1150_up", this);
    pf_vf_mux_scbd_1151_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1151_up", this);
    pf_vf_mux_scbd_1152_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1152_up", this);
    pf_vf_mux_scbd_1153_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1153_up", this);
    pf_vf_mux_scbd_1154_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1154_up", this);
    pf_vf_mux_scbd_1155_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1155_up", this);
    pf_vf_mux_scbd_1156_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1156_up", this);
    pf_vf_mux_scbd_1157_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1157_up", this);
    pf_vf_mux_scbd_1158_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1158_up", this);
    pf_vf_mux_scbd_1159_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1159_up", this);
    pf_vf_mux_scbd_1160_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1160_up", this);
    pf_vf_mux_scbd_1161_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1161_up", this);
    pf_vf_mux_scbd_1162_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1162_up", this);
    pf_vf_mux_scbd_1163_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1163_up", this);
    pf_vf_mux_scbd_1164_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1164_up", this);
    pf_vf_mux_scbd_1165_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1165_up", this);
    pf_vf_mux_scbd_1166_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1166_up", this);
    pf_vf_mux_scbd_1167_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1167_up", this);
    pf_vf_mux_scbd_1168_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1168_up", this);
    pf_vf_mux_scbd_1169_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1169_up", this);
    pf_vf_mux_scbd_1170_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1170_up", this);
    pf_vf_mux_scbd_1171_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1171_up", this);
    pf_vf_mux_scbd_1172_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1172_up", this);
    pf_vf_mux_scbd_1173_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1173_up", this);
    pf_vf_mux_scbd_1174_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1174_up", this);
    pf_vf_mux_scbd_1175_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1175_up", this);
    pf_vf_mux_scbd_1176_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1176_up", this);
    pf_vf_mux_scbd_1177_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1177_up", this);
    pf_vf_mux_scbd_1178_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1178_up", this);
    pf_vf_mux_scbd_1179_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1179_up", this);
    pf_vf_mux_scbd_1180_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1180_up", this);
    pf_vf_mux_scbd_1181_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1181_up", this);
    pf_vf_mux_scbd_1182_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1182_up", this);
    pf_vf_mux_scbd_1183_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1183_up", this);
    pf_vf_mux_scbd_1184_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1184_up", this);
    pf_vf_mux_scbd_1185_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1185_up", this);
    pf_vf_mux_scbd_1186_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1186_up", this);
    pf_vf_mux_scbd_1187_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1187_up", this);
    pf_vf_mux_scbd_1188_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1188_up", this);
    pf_vf_mux_scbd_1189_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1189_up", this);
    pf_vf_mux_scbd_1190_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1190_up", this);
    pf_vf_mux_scbd_1191_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1191_up", this);
    pf_vf_mux_scbd_1192_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1192_up", this);
    pf_vf_mux_scbd_1193_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1193_up", this);
    pf_vf_mux_scbd_1194_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1194_up", this);
    pf_vf_mux_scbd_1195_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1195_up", this);
    pf_vf_mux_scbd_1196_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1196_up", this);
    pf_vf_mux_scbd_1197_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1197_up", this);
    pf_vf_mux_scbd_1198_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1198_up", this);
    pf_vf_mux_scbd_1199_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1199_up", this);
    pf_vf_mux_scbd_1200_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1200_up", this);
    pf_vf_mux_scbd_1201_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1201_up", this);
    pf_vf_mux_scbd_1202_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1202_up", this);
    pf_vf_mux_scbd_1203_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1203_up", this);
    pf_vf_mux_scbd_1204_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1204_up", this);
    pf_vf_mux_scbd_1205_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1205_up", this);
    pf_vf_mux_scbd_1206_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1206_up", this);
    pf_vf_mux_scbd_1207_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1207_up", this);
    pf_vf_mux_scbd_1208_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1208_up", this);
    pf_vf_mux_scbd_1209_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1209_up", this);
    pf_vf_mux_scbd_1210_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1210_up", this);
    pf_vf_mux_scbd_1211_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1211_up", this);
    pf_vf_mux_scbd_1212_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1212_up", this);
    pf_vf_mux_scbd_1213_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1213_up", this);
    pf_vf_mux_scbd_1214_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1214_up", this);
    pf_vf_mux_scbd_1215_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1215_up", this);
    pf_vf_mux_scbd_1216_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1216_up", this);
    pf_vf_mux_scbd_1217_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1217_up", this);
    pf_vf_mux_scbd_1218_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1218_up", this);
    pf_vf_mux_scbd_1219_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1219_up", this);
    pf_vf_mux_scbd_1220_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1220_up", this);
    pf_vf_mux_scbd_1221_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1221_up", this);
    pf_vf_mux_scbd_1222_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1222_up", this);
    pf_vf_mux_scbd_1223_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1223_up", this);
    pf_vf_mux_scbd_1224_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1224_up", this);
    pf_vf_mux_scbd_1225_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1225_up", this);
    pf_vf_mux_scbd_1226_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1226_up", this);
    pf_vf_mux_scbd_1227_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1227_up", this);
    pf_vf_mux_scbd_1228_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1228_up", this);
    pf_vf_mux_scbd_1229_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1229_up", this);
    pf_vf_mux_scbd_1230_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1230_up", this);
    pf_vf_mux_scbd_1231_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1231_up", this);
    pf_vf_mux_scbd_1232_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1232_up", this);
    pf_vf_mux_scbd_1233_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1233_up", this);
    pf_vf_mux_scbd_1234_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1234_up", this);
    pf_vf_mux_scbd_1235_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1235_up", this);
    pf_vf_mux_scbd_1236_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1236_up", this);
    pf_vf_mux_scbd_1237_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1237_up", this);
    pf_vf_mux_scbd_1238_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1238_up", this);
    pf_vf_mux_scbd_1239_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1239_up", this);
    pf_vf_mux_scbd_1240_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1240_up", this);
    pf_vf_mux_scbd_1241_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1241_up", this);
    pf_vf_mux_scbd_1242_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1242_up", this);
    pf_vf_mux_scbd_1243_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1243_up", this);
    pf_vf_mux_scbd_1244_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1244_up", this);
    pf_vf_mux_scbd_1245_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1245_up", this);
    pf_vf_mux_scbd_1246_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1246_up", this);
    pf_vf_mux_scbd_1247_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1247_up", this);
    pf_vf_mux_scbd_1248_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1248_up", this);
    pf_vf_mux_scbd_1249_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1249_up", this);
    pf_vf_mux_scbd_1250_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1250_up", this);
    pf_vf_mux_scbd_1251_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1251_up", this);
    pf_vf_mux_scbd_1252_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1252_up", this);
    pf_vf_mux_scbd_1253_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1253_up", this);
    pf_vf_mux_scbd_1254_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1254_up", this);
    pf_vf_mux_scbd_1255_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1255_up", this);
    pf_vf_mux_scbd_1256_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1256_up", this);
    pf_vf_mux_scbd_1257_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1257_up", this);
    pf_vf_mux_scbd_1258_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1258_up", this);
    pf_vf_mux_scbd_1259_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1259_up", this);
    pf_vf_mux_scbd_1260_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1260_up", this);
    pf_vf_mux_scbd_1261_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1261_up", this);
    pf_vf_mux_scbd_1262_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1262_up", this);
    pf_vf_mux_scbd_1263_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1263_up", this);
    pf_vf_mux_scbd_1264_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1264_up", this);
    pf_vf_mux_scbd_1265_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1265_up", this);
    pf_vf_mux_scbd_1266_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1266_up", this);
    pf_vf_mux_scbd_1267_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1267_up", this);
    pf_vf_mux_scbd_1268_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1268_up", this);
    pf_vf_mux_scbd_1269_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1269_up", this);
    pf_vf_mux_scbd_1270_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1270_up", this);
    pf_vf_mux_scbd_1271_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1271_up", this);
    pf_vf_mux_scbd_1272_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1272_up", this);
    pf_vf_mux_scbd_1273_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1273_up", this);
    pf_vf_mux_scbd_1274_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1274_up", this);
    pf_vf_mux_scbd_1275_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1275_up", this);
    pf_vf_mux_scbd_1276_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1276_up", this);
    pf_vf_mux_scbd_1277_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1277_up", this);
    pf_vf_mux_scbd_1278_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1278_up", this);
    pf_vf_mux_scbd_1279_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1279_up", this);
    pf_vf_mux_scbd_1280_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1280_up", this);
    pf_vf_mux_scbd_1281_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1281_up", this);
    pf_vf_mux_scbd_1282_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1282_up", this);
    pf_vf_mux_scbd_1283_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1283_up", this);
    pf_vf_mux_scbd_1284_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1284_up", this);
    pf_vf_mux_scbd_1285_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1285_up", this);
    pf_vf_mux_scbd_1286_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1286_up", this);
    pf_vf_mux_scbd_1287_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1287_up", this);
    pf_vf_mux_scbd_1288_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1288_up", this);
    pf_vf_mux_scbd_1289_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1289_up", this);
    pf_vf_mux_scbd_1290_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1290_up", this);
    pf_vf_mux_scbd_1291_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1291_up", this);
    pf_vf_mux_scbd_1292_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1292_up", this);
    pf_vf_mux_scbd_1293_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1293_up", this);
    pf_vf_mux_scbd_1294_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1294_up", this);
    pf_vf_mux_scbd_1295_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1295_up", this);
    pf_vf_mux_scbd_1296_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1296_up", this);
    pf_vf_mux_scbd_1297_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1297_up", this);
    pf_vf_mux_scbd_1298_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1298_up", this);
    pf_vf_mux_scbd_1299_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1299_up", this);
    pf_vf_mux_scbd_1300_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1300_up", this);
    pf_vf_mux_scbd_1301_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1301_up", this);
    pf_vf_mux_scbd_1302_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1302_up", this);
    pf_vf_mux_scbd_1303_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1303_up", this);
    pf_vf_mux_scbd_1304_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1304_up", this);
    pf_vf_mux_scbd_1305_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1305_up", this);
    pf_vf_mux_scbd_1306_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1306_up", this);
    pf_vf_mux_scbd_1307_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1307_up", this);
    pf_vf_mux_scbd_1308_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1308_up", this);
    pf_vf_mux_scbd_1309_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1309_up", this);
    pf_vf_mux_scbd_1310_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1310_up", this);
    pf_vf_mux_scbd_1311_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1311_up", this);
    pf_vf_mux_scbd_1312_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1312_up", this);
    pf_vf_mux_scbd_1313_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1313_up", this);
    pf_vf_mux_scbd_1314_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1314_up", this);
    pf_vf_mux_scbd_1315_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1315_up", this);
    pf_vf_mux_scbd_1316_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1316_up", this);
    pf_vf_mux_scbd_1317_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1317_up", this);
    pf_vf_mux_scbd_1318_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1318_up", this);
    pf_vf_mux_scbd_1319_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1319_up", this);
    pf_vf_mux_scbd_1320_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1320_up", this);
    pf_vf_mux_scbd_1321_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1321_up", this);
    pf_vf_mux_scbd_1322_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1322_up", this);
    pf_vf_mux_scbd_1323_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1323_up", this);
    pf_vf_mux_scbd_1324_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1324_up", this);
    pf_vf_mux_scbd_1325_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1325_up", this);
    pf_vf_mux_scbd_1326_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1326_up", this);
    pf_vf_mux_scbd_1327_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1327_up", this);
    pf_vf_mux_scbd_1328_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1328_up", this);
    pf_vf_mux_scbd_1329_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1329_up", this);
    pf_vf_mux_scbd_1330_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1330_up", this);
    pf_vf_mux_scbd_1331_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1331_up", this);
    pf_vf_mux_scbd_1332_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1332_up", this);
    pf_vf_mux_scbd_1333_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1333_up", this);
    pf_vf_mux_scbd_1334_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1334_up", this);
    pf_vf_mux_scbd_1335_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1335_up", this);
    pf_vf_mux_scbd_1336_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1336_up", this);
    pf_vf_mux_scbd_1337_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1337_up", this);
    pf_vf_mux_scbd_1338_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1338_up", this);
    pf_vf_mux_scbd_1339_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1339_up", this);
    pf_vf_mux_scbd_1340_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1340_up", this);
    pf_vf_mux_scbd_1341_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1341_up", this);
    pf_vf_mux_scbd_1342_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1342_up", this);
    pf_vf_mux_scbd_1343_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1343_up", this);
    pf_vf_mux_scbd_1344_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1344_up", this);
    pf_vf_mux_scbd_1345_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1345_up", this);
    pf_vf_mux_scbd_1346_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1346_up", this);
    pf_vf_mux_scbd_1347_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1347_up", this);
    pf_vf_mux_scbd_1348_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1348_up", this);
    pf_vf_mux_scbd_1349_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1349_up", this);
    pf_vf_mux_scbd_1350_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1350_up", this);
    pf_vf_mux_scbd_1351_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1351_up", this);
    pf_vf_mux_scbd_1352_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1352_up", this);
    pf_vf_mux_scbd_1353_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1353_up", this);
    pf_vf_mux_scbd_1354_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1354_up", this);
    pf_vf_mux_scbd_1355_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1355_up", this);
    pf_vf_mux_scbd_1356_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1356_up", this);
    pf_vf_mux_scbd_1357_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1357_up", this);
    pf_vf_mux_scbd_1358_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1358_up", this);
    pf_vf_mux_scbd_1359_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1359_up", this);
    pf_vf_mux_scbd_1360_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1360_up", this);
    pf_vf_mux_scbd_1361_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1361_up", this);
    pf_vf_mux_scbd_1362_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1362_up", this);
    pf_vf_mux_scbd_1363_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1363_up", this);
    pf_vf_mux_scbd_1364_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1364_up", this);
    pf_vf_mux_scbd_1365_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1365_up", this);
    pf_vf_mux_scbd_1366_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1366_up", this);
    pf_vf_mux_scbd_1367_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1367_up", this);
    pf_vf_mux_scbd_1368_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1368_up", this);
    pf_vf_mux_scbd_1369_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1369_up", this);
    pf_vf_mux_scbd_1370_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1370_up", this);
    pf_vf_mux_scbd_1371_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1371_up", this);
    pf_vf_mux_scbd_1372_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1372_up", this);
    pf_vf_mux_scbd_1373_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1373_up", this);
    pf_vf_mux_scbd_1374_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1374_up", this);
    pf_vf_mux_scbd_1375_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1375_up", this);
    pf_vf_mux_scbd_1376_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1376_up", this);
    pf_vf_mux_scbd_1377_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1377_up", this);
    pf_vf_mux_scbd_1378_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1378_up", this);
    pf_vf_mux_scbd_1379_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1379_up", this);
    pf_vf_mux_scbd_1380_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1380_up", this);
    pf_vf_mux_scbd_1381_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1381_up", this);
    pf_vf_mux_scbd_1382_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1382_up", this);
    pf_vf_mux_scbd_1383_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1383_up", this);
    pf_vf_mux_scbd_1384_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1384_up", this);
    pf_vf_mux_scbd_1385_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1385_up", this);
    pf_vf_mux_scbd_1386_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1386_up", this);
    pf_vf_mux_scbd_1387_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1387_up", this);
    pf_vf_mux_scbd_1388_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1388_up", this);
    pf_vf_mux_scbd_1389_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1389_up", this);
    pf_vf_mux_scbd_1390_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1390_up", this);
    pf_vf_mux_scbd_1391_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1391_up", this);
    pf_vf_mux_scbd_1392_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1392_up", this);
    pf_vf_mux_scbd_1393_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1393_up", this);
    pf_vf_mux_scbd_1394_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1394_up", this);
    pf_vf_mux_scbd_1395_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1395_up", this);
    pf_vf_mux_scbd_1396_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1396_up", this);
    pf_vf_mux_scbd_1397_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1397_up", this);
    pf_vf_mux_scbd_1398_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1398_up", this);
    pf_vf_mux_scbd_1399_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1399_up", this);
    pf_vf_mux_scbd_1400_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1400_up", this);
    pf_vf_mux_scbd_1401_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1401_up", this);
    pf_vf_mux_scbd_1402_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1402_up", this);
    pf_vf_mux_scbd_1403_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1403_up", this);
    pf_vf_mux_scbd_1404_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1404_up", this);
    pf_vf_mux_scbd_1405_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1405_up", this);
    pf_vf_mux_scbd_1406_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1406_up", this);
    pf_vf_mux_scbd_1407_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1407_up", this);
    pf_vf_mux_scbd_1408_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1408_up", this);
    pf_vf_mux_scbd_1409_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1409_up", this);
    pf_vf_mux_scbd_1410_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1410_up", this);
    pf_vf_mux_scbd_1411_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1411_up", this);
    pf_vf_mux_scbd_1412_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1412_up", this);
    pf_vf_mux_scbd_1413_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1413_up", this);
    pf_vf_mux_scbd_1414_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1414_up", this);
    pf_vf_mux_scbd_1415_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1415_up", this);
    pf_vf_mux_scbd_1416_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1416_up", this);
    pf_vf_mux_scbd_1417_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1417_up", this);
    pf_vf_mux_scbd_1418_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1418_up", this);
    pf_vf_mux_scbd_1419_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1419_up", this);
    pf_vf_mux_scbd_1420_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1420_up", this);
    pf_vf_mux_scbd_1421_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1421_up", this);
    pf_vf_mux_scbd_1422_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1422_up", this);
    pf_vf_mux_scbd_1423_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1423_up", this);
    pf_vf_mux_scbd_1424_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1424_up", this);
    pf_vf_mux_scbd_1425_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1425_up", this);
    pf_vf_mux_scbd_1426_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1426_up", this);
    pf_vf_mux_scbd_1427_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1427_up", this);
    pf_vf_mux_scbd_1428_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1428_up", this);
    pf_vf_mux_scbd_1429_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1429_up", this);
    pf_vf_mux_scbd_1430_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1430_up", this);
    pf_vf_mux_scbd_1431_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1431_up", this);
    pf_vf_mux_scbd_1432_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1432_up", this);
    pf_vf_mux_scbd_1433_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1433_up", this);
    pf_vf_mux_scbd_1434_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1434_up", this);
    pf_vf_mux_scbd_1435_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1435_up", this);
    pf_vf_mux_scbd_1436_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1436_up", this);
    pf_vf_mux_scbd_1437_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1437_up", this);
    pf_vf_mux_scbd_1438_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1438_up", this);
    pf_vf_mux_scbd_1439_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1439_up", this);
    pf_vf_mux_scbd_1440_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1440_up", this);
    pf_vf_mux_scbd_1441_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1441_up", this);
    pf_vf_mux_scbd_1442_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1442_up", this);
    pf_vf_mux_scbd_1443_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1443_up", this);
    pf_vf_mux_scbd_1444_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1444_up", this);
    pf_vf_mux_scbd_1445_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1445_up", this);
    pf_vf_mux_scbd_1446_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1446_up", this);
    pf_vf_mux_scbd_1447_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1447_up", this);
    pf_vf_mux_scbd_1448_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1448_up", this);
    pf_vf_mux_scbd_1449_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1449_up", this);
    pf_vf_mux_scbd_1450_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1450_up", this);
    pf_vf_mux_scbd_1451_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1451_up", this);
    pf_vf_mux_scbd_1452_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1452_up", this);
    pf_vf_mux_scbd_1453_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1453_up", this);
    pf_vf_mux_scbd_1454_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1454_up", this);
    pf_vf_mux_scbd_1455_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1455_up", this);
    pf_vf_mux_scbd_1456_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1456_up", this);
    pf_vf_mux_scbd_1457_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1457_up", this);
    pf_vf_mux_scbd_1458_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1458_up", this);
    pf_vf_mux_scbd_1459_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1459_up", this);
    pf_vf_mux_scbd_1460_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1460_up", this);
    pf_vf_mux_scbd_1461_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1461_up", this);
    pf_vf_mux_scbd_1462_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1462_up", this);
    pf_vf_mux_scbd_1463_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1463_up", this);
    pf_vf_mux_scbd_1464_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1464_up", this);
    pf_vf_mux_scbd_1465_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1465_up", this);
    pf_vf_mux_scbd_1466_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1466_up", this);
    pf_vf_mux_scbd_1467_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1467_up", this);
    pf_vf_mux_scbd_1468_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1468_up", this);
    pf_vf_mux_scbd_1469_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1469_up", this);
    pf_vf_mux_scbd_1470_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1470_up", this);
    pf_vf_mux_scbd_1471_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1471_up", this);
    pf_vf_mux_scbd_1472_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1472_up", this);
    pf_vf_mux_scbd_1473_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1473_up", this);
    pf_vf_mux_scbd_1474_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1474_up", this);
    pf_vf_mux_scbd_1475_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1475_up", this);
    pf_vf_mux_scbd_1476_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1476_up", this);
    pf_vf_mux_scbd_1477_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1477_up", this);
    pf_vf_mux_scbd_1478_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1478_up", this);
    pf_vf_mux_scbd_1479_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1479_up", this);
    pf_vf_mux_scbd_1480_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1480_up", this);
    pf_vf_mux_scbd_1481_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1481_up", this);
    pf_vf_mux_scbd_1482_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1482_up", this);
    pf_vf_mux_scbd_1483_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1483_up", this);
    pf_vf_mux_scbd_1484_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1484_up", this);
    pf_vf_mux_scbd_1485_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1485_up", this);
    pf_vf_mux_scbd_1486_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1486_up", this);
    pf_vf_mux_scbd_1487_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1487_up", this);
    pf_vf_mux_scbd_1488_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1488_up", this);
    pf_vf_mux_scbd_1489_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1489_up", this);
    pf_vf_mux_scbd_1490_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1490_up", this);
    pf_vf_mux_scbd_1491_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1491_up", this);
    pf_vf_mux_scbd_1492_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1492_up", this);
    pf_vf_mux_scbd_1493_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1493_up", this);
    pf_vf_mux_scbd_1494_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1494_up", this);
    pf_vf_mux_scbd_1495_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1495_up", this);
    pf_vf_mux_scbd_1496_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1496_up", this);
    pf_vf_mux_scbd_1497_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1497_up", this);
    pf_vf_mux_scbd_1498_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1498_up", this);
    pf_vf_mux_scbd_1499_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1499_up", this);
    pf_vf_mux_scbd_1500_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1500_up", this);
    pf_vf_mux_scbd_1501_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1501_up", this);
    pf_vf_mux_scbd_1502_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1502_up", this);
    pf_vf_mux_scbd_1503_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1503_up", this);
    pf_vf_mux_scbd_1504_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1504_up", this);
    pf_vf_mux_scbd_1505_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1505_up", this);
    pf_vf_mux_scbd_1506_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1506_up", this);
    pf_vf_mux_scbd_1507_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1507_up", this);
    pf_vf_mux_scbd_1508_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1508_up", this);
    pf_vf_mux_scbd_1509_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1509_up", this);
    pf_vf_mux_scbd_1510_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1510_up", this);
    pf_vf_mux_scbd_1511_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1511_up", this);
    pf_vf_mux_scbd_1512_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1512_up", this);
    pf_vf_mux_scbd_1513_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1513_up", this);
    pf_vf_mux_scbd_1514_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1514_up", this);
    pf_vf_mux_scbd_1515_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1515_up", this);
    pf_vf_mux_scbd_1516_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1516_up", this);
    pf_vf_mux_scbd_1517_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1517_up", this);
    pf_vf_mux_scbd_1518_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1518_up", this);
    pf_vf_mux_scbd_1519_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1519_up", this);
    pf_vf_mux_scbd_1520_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1520_up", this);
    pf_vf_mux_scbd_1521_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1521_up", this);
    pf_vf_mux_scbd_1522_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1522_up", this);
    pf_vf_mux_scbd_1523_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1523_up", this);
    pf_vf_mux_scbd_1524_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1524_up", this);
    pf_vf_mux_scbd_1525_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1525_up", this);
    pf_vf_mux_scbd_1526_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1526_up", this);
    pf_vf_mux_scbd_1527_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1527_up", this);
    pf_vf_mux_scbd_1528_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1528_up", this);
    pf_vf_mux_scbd_1529_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1529_up", this);
    pf_vf_mux_scbd_1530_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1530_up", this);
    pf_vf_mux_scbd_1531_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1531_up", this);
    pf_vf_mux_scbd_1532_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1532_up", this);
    pf_vf_mux_scbd_1533_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1533_up", this);
    pf_vf_mux_scbd_1534_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1534_up", this);
    pf_vf_mux_scbd_1535_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1535_up", this);
    pf_vf_mux_scbd_1536_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1536_up", this);
    pf_vf_mux_scbd_1537_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1537_up", this);
    pf_vf_mux_scbd_1538_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1538_up", this);
    pf_vf_mux_scbd_1539_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1539_up", this);
    pf_vf_mux_scbd_1540_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1540_up", this);
    pf_vf_mux_scbd_1541_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1541_up", this);
    pf_vf_mux_scbd_1542_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1542_up", this);
    pf_vf_mux_scbd_1543_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1543_up", this);
    pf_vf_mux_scbd_1544_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1544_up", this);
    pf_vf_mux_scbd_1545_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1545_up", this);
    pf_vf_mux_scbd_1546_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1546_up", this);
    pf_vf_mux_scbd_1547_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1547_up", this);
    pf_vf_mux_scbd_1548_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1548_up", this);
    pf_vf_mux_scbd_1549_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1549_up", this);
    pf_vf_mux_scbd_1550_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1550_up", this);
    pf_vf_mux_scbd_1551_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1551_up", this);
    pf_vf_mux_scbd_1552_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1552_up", this);
    pf_vf_mux_scbd_1553_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1553_up", this);
    pf_vf_mux_scbd_1554_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1554_up", this);
    pf_vf_mux_scbd_1555_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1555_up", this);
    pf_vf_mux_scbd_1556_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1556_up", this);
    pf_vf_mux_scbd_1557_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1557_up", this);
    pf_vf_mux_scbd_1558_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1558_up", this);
    pf_vf_mux_scbd_1559_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1559_up", this);
    pf_vf_mux_scbd_1560_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1560_up", this);
    pf_vf_mux_scbd_1561_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1561_up", this);
    pf_vf_mux_scbd_1562_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1562_up", this);
    pf_vf_mux_scbd_1563_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1563_up", this);
    pf_vf_mux_scbd_1564_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1564_up", this);
    pf_vf_mux_scbd_1565_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1565_up", this);
    pf_vf_mux_scbd_1566_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1566_up", this);
    pf_vf_mux_scbd_1567_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1567_up", this);
    pf_vf_mux_scbd_1568_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1568_up", this);
    pf_vf_mux_scbd_1569_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1569_up", this);
    pf_vf_mux_scbd_1570_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1570_up", this);
    pf_vf_mux_scbd_1571_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1571_up", this);
    pf_vf_mux_scbd_1572_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1572_up", this);
    pf_vf_mux_scbd_1573_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1573_up", this);
    pf_vf_mux_scbd_1574_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1574_up", this);
    pf_vf_mux_scbd_1575_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1575_up", this);
    pf_vf_mux_scbd_1576_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1576_up", this);
    pf_vf_mux_scbd_1577_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1577_up", this);
    pf_vf_mux_scbd_1578_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1578_up", this);
    pf_vf_mux_scbd_1579_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1579_up", this);
    pf_vf_mux_scbd_1580_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1580_up", this);
    pf_vf_mux_scbd_1581_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1581_up", this);
    pf_vf_mux_scbd_1582_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1582_up", this);
    pf_vf_mux_scbd_1583_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1583_up", this);
    pf_vf_mux_scbd_1584_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1584_up", this);
    pf_vf_mux_scbd_1585_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1585_up", this);
    pf_vf_mux_scbd_1586_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1586_up", this);
    pf_vf_mux_scbd_1587_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1587_up", this);
    pf_vf_mux_scbd_1588_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1588_up", this);
    pf_vf_mux_scbd_1589_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1589_up", this);
    pf_vf_mux_scbd_1590_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1590_up", this);
    pf_vf_mux_scbd_1591_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1591_up", this);
    pf_vf_mux_scbd_1592_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1592_up", this);
    pf_vf_mux_scbd_1593_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1593_up", this);
    pf_vf_mux_scbd_1594_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1594_up", this);
    pf_vf_mux_scbd_1595_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1595_up", this);
    pf_vf_mux_scbd_1596_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1596_up", this);
    pf_vf_mux_scbd_1597_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1597_up", this);
    pf_vf_mux_scbd_1598_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1598_up", this);
    pf_vf_mux_scbd_1599_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1599_up", this);
    pf_vf_mux_scbd_1600_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1600_up", this);
    pf_vf_mux_scbd_1601_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1601_up", this);
    pf_vf_mux_scbd_1602_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1602_up", this);
    pf_vf_mux_scbd_1603_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1603_up", this);
    pf_vf_mux_scbd_1604_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1604_up", this);
    pf_vf_mux_scbd_1605_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1605_up", this);
    pf_vf_mux_scbd_1606_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1606_up", this);
    pf_vf_mux_scbd_1607_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1607_up", this);
    pf_vf_mux_scbd_1608_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1608_up", this);
    pf_vf_mux_scbd_1609_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1609_up", this);
    pf_vf_mux_scbd_1610_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1610_up", this);
    pf_vf_mux_scbd_1611_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1611_up", this);
    pf_vf_mux_scbd_1612_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1612_up", this);
    pf_vf_mux_scbd_1613_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1613_up", this);
    pf_vf_mux_scbd_1614_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1614_up", this);
    pf_vf_mux_scbd_1615_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1615_up", this);
    pf_vf_mux_scbd_1616_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1616_up", this);
    pf_vf_mux_scbd_1617_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1617_up", this);
    pf_vf_mux_scbd_1618_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1618_up", this);
    pf_vf_mux_scbd_1619_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1619_up", this);
    pf_vf_mux_scbd_1620_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1620_up", this);
    pf_vf_mux_scbd_1621_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1621_up", this);
    pf_vf_mux_scbd_1622_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1622_up", this);
    pf_vf_mux_scbd_1623_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1623_up", this);
    pf_vf_mux_scbd_1624_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1624_up", this);
    pf_vf_mux_scbd_1625_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1625_up", this);
    pf_vf_mux_scbd_1626_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1626_up", this);
    pf_vf_mux_scbd_1627_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1627_up", this);
    pf_vf_mux_scbd_1628_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1628_up", this);
    pf_vf_mux_scbd_1629_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1629_up", this);
    pf_vf_mux_scbd_1630_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1630_up", this);
    pf_vf_mux_scbd_1631_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1631_up", this);
    pf_vf_mux_scbd_1632_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1632_up", this);
    pf_vf_mux_scbd_1633_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1633_up", this);
    pf_vf_mux_scbd_1634_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1634_up", this);
    pf_vf_mux_scbd_1635_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1635_up", this);
    pf_vf_mux_scbd_1636_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1636_up", this);
    pf_vf_mux_scbd_1637_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1637_up", this);
    pf_vf_mux_scbd_1638_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1638_up", this);
    pf_vf_mux_scbd_1639_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1639_up", this);
    pf_vf_mux_scbd_1640_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1640_up", this);
    pf_vf_mux_scbd_1641_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1641_up", this);
    pf_vf_mux_scbd_1642_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1642_up", this);
    pf_vf_mux_scbd_1643_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1643_up", this);
    pf_vf_mux_scbd_1644_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1644_up", this);
    pf_vf_mux_scbd_1645_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1645_up", this);
    pf_vf_mux_scbd_1646_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1646_up", this);
    pf_vf_mux_scbd_1647_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1647_up", this);
    pf_vf_mux_scbd_1648_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1648_up", this);
    pf_vf_mux_scbd_1649_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1649_up", this);
    pf_vf_mux_scbd_1650_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1650_up", this);
    pf_vf_mux_scbd_1651_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1651_up", this);
    pf_vf_mux_scbd_1652_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1652_up", this);
    pf_vf_mux_scbd_1653_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1653_up", this);
    pf_vf_mux_scbd_1654_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1654_up", this);
    pf_vf_mux_scbd_1655_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1655_up", this);
    pf_vf_mux_scbd_1656_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1656_up", this);
    pf_vf_mux_scbd_1657_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1657_up", this);
    pf_vf_mux_scbd_1658_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1658_up", this);
    pf_vf_mux_scbd_1659_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1659_up", this);
    pf_vf_mux_scbd_1660_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1660_up", this);
    pf_vf_mux_scbd_1661_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1661_up", this);
    pf_vf_mux_scbd_1662_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1662_up", this);
    pf_vf_mux_scbd_1663_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1663_up", this);
    pf_vf_mux_scbd_1664_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1664_up", this);
    pf_vf_mux_scbd_1665_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1665_up", this);
    pf_vf_mux_scbd_1666_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1666_up", this);
    pf_vf_mux_scbd_1667_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1667_up", this);
    pf_vf_mux_scbd_1668_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1668_up", this);
    pf_vf_mux_scbd_1669_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1669_up", this);
    pf_vf_mux_scbd_1670_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1670_up", this);
    pf_vf_mux_scbd_1671_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1671_up", this);
    pf_vf_mux_scbd_1672_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1672_up", this);
    pf_vf_mux_scbd_1673_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1673_up", this);
    pf_vf_mux_scbd_1674_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1674_up", this);
    pf_vf_mux_scbd_1675_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1675_up", this);
    pf_vf_mux_scbd_1676_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1676_up", this);
    pf_vf_mux_scbd_1677_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1677_up", this);
    pf_vf_mux_scbd_1678_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1678_up", this);
    pf_vf_mux_scbd_1679_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1679_up", this);
    pf_vf_mux_scbd_1680_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1680_up", this);
    pf_vf_mux_scbd_1681_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1681_up", this);
    pf_vf_mux_scbd_1682_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1682_up", this);
    pf_vf_mux_scbd_1683_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1683_up", this);
    pf_vf_mux_scbd_1684_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1684_up", this);
    pf_vf_mux_scbd_1685_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1685_up", this);
    pf_vf_mux_scbd_1686_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1686_up", this);
    pf_vf_mux_scbd_1687_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1687_up", this);
    pf_vf_mux_scbd_1688_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1688_up", this);
    pf_vf_mux_scbd_1689_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1689_up", this);
    pf_vf_mux_scbd_1690_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1690_up", this);
    pf_vf_mux_scbd_1691_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1691_up", this);
    pf_vf_mux_scbd_1692_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1692_up", this);
    pf_vf_mux_scbd_1693_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1693_up", this);
    pf_vf_mux_scbd_1694_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1694_up", this);
    pf_vf_mux_scbd_1695_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1695_up", this);
    pf_vf_mux_scbd_1696_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1696_up", this);
    pf_vf_mux_scbd_1697_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1697_up", this);
    pf_vf_mux_scbd_1698_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1698_up", this);
    pf_vf_mux_scbd_1699_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1699_up", this);
    pf_vf_mux_scbd_1700_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1700_up", this);
    pf_vf_mux_scbd_1701_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1701_up", this);
    pf_vf_mux_scbd_1702_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1702_up", this);
    pf_vf_mux_scbd_1703_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1703_up", this);
    pf_vf_mux_scbd_1704_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1704_up", this);
    pf_vf_mux_scbd_1705_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1705_up", this);
    pf_vf_mux_scbd_1706_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1706_up", this);
    pf_vf_mux_scbd_1707_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1707_up", this);
    pf_vf_mux_scbd_1708_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1708_up", this);
    pf_vf_mux_scbd_1709_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1709_up", this);
    pf_vf_mux_scbd_1710_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1710_up", this);
    pf_vf_mux_scbd_1711_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1711_up", this);
    pf_vf_mux_scbd_1712_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1712_up", this);
    pf_vf_mux_scbd_1713_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1713_up", this);
    pf_vf_mux_scbd_1714_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1714_up", this);
    pf_vf_mux_scbd_1715_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1715_up", this);
    pf_vf_mux_scbd_1716_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1716_up", this);
    pf_vf_mux_scbd_1717_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1717_up", this);
    pf_vf_mux_scbd_1718_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1718_up", this);
    pf_vf_mux_scbd_1719_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1719_up", this);
    pf_vf_mux_scbd_1720_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1720_up", this);
    pf_vf_mux_scbd_1721_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1721_up", this);
    pf_vf_mux_scbd_1722_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1722_up", this);
    pf_vf_mux_scbd_1723_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1723_up", this);
    pf_vf_mux_scbd_1724_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1724_up", this);
    pf_vf_mux_scbd_1725_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1725_up", this);
    pf_vf_mux_scbd_1726_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1726_up", this);
    pf_vf_mux_scbd_1727_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1727_up", this);
    pf_vf_mux_scbd_1728_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1728_up", this);
    pf_vf_mux_scbd_1729_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1729_up", this);
    pf_vf_mux_scbd_1730_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1730_up", this);
    pf_vf_mux_scbd_1731_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1731_up", this);
    pf_vf_mux_scbd_1732_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1732_up", this);
    pf_vf_mux_scbd_1733_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1733_up", this);
    pf_vf_mux_scbd_1734_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1734_up", this);
    pf_vf_mux_scbd_1735_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1735_up", this);
    pf_vf_mux_scbd_1736_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1736_up", this);
    pf_vf_mux_scbd_1737_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1737_up", this);
    pf_vf_mux_scbd_1738_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1738_up", this);
    pf_vf_mux_scbd_1739_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1739_up", this);
    pf_vf_mux_scbd_1740_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1740_up", this);
    pf_vf_mux_scbd_1741_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1741_up", this);
    pf_vf_mux_scbd_1742_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1742_up", this);
    pf_vf_mux_scbd_1743_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1743_up", this);
    pf_vf_mux_scbd_1744_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1744_up", this);
    pf_vf_mux_scbd_1745_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1745_up", this);
    pf_vf_mux_scbd_1746_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1746_up", this);
    pf_vf_mux_scbd_1747_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1747_up", this);
    pf_vf_mux_scbd_1748_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1748_up", this);
    pf_vf_mux_scbd_1749_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1749_up", this);
    pf_vf_mux_scbd_1750_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1750_up", this);
    pf_vf_mux_scbd_1751_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1751_up", this);
    pf_vf_mux_scbd_1752_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1752_up", this);
    pf_vf_mux_scbd_1753_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1753_up", this);
    pf_vf_mux_scbd_1754_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1754_up", this);
    pf_vf_mux_scbd_1755_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1755_up", this);
    pf_vf_mux_scbd_1756_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1756_up", this);
    pf_vf_mux_scbd_1757_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1757_up", this);
    pf_vf_mux_scbd_1758_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1758_up", this);
    pf_vf_mux_scbd_1759_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1759_up", this);
    pf_vf_mux_scbd_1760_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1760_up", this);
    pf_vf_mux_scbd_1761_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1761_up", this);
    pf_vf_mux_scbd_1762_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1762_up", this);
    pf_vf_mux_scbd_1763_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1763_up", this);
    pf_vf_mux_scbd_1764_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1764_up", this);
    pf_vf_mux_scbd_1765_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1765_up", this);
    pf_vf_mux_scbd_1766_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1766_up", this);
    pf_vf_mux_scbd_1767_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1767_up", this);
    pf_vf_mux_scbd_1768_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1768_up", this);
    pf_vf_mux_scbd_1769_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1769_up", this);
    pf_vf_mux_scbd_1770_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1770_up", this);
    pf_vf_mux_scbd_1771_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1771_up", this);
    pf_vf_mux_scbd_1772_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1772_up", this);
    pf_vf_mux_scbd_1773_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1773_up", this);
    pf_vf_mux_scbd_1774_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1774_up", this);
    pf_vf_mux_scbd_1775_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1775_up", this);
    pf_vf_mux_scbd_1776_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1776_up", this);
    pf_vf_mux_scbd_1777_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1777_up", this);
    pf_vf_mux_scbd_1778_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1778_up", this);
    pf_vf_mux_scbd_1779_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1779_up", this);
    pf_vf_mux_scbd_1780_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1780_up", this);
    pf_vf_mux_scbd_1781_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1781_up", this);
    pf_vf_mux_scbd_1782_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1782_up", this);
    pf_vf_mux_scbd_1783_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1783_up", this);
    pf_vf_mux_scbd_1784_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1784_up", this);
    pf_vf_mux_scbd_1785_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1785_up", this);
    pf_vf_mux_scbd_1786_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1786_up", this);
    pf_vf_mux_scbd_1787_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1787_up", this);
    pf_vf_mux_scbd_1788_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1788_up", this);
    pf_vf_mux_scbd_1789_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1789_up", this);
    pf_vf_mux_scbd_1790_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1790_up", this);
    pf_vf_mux_scbd_1791_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1791_up", this);
    pf_vf_mux_scbd_1792_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1792_up", this);
    pf_vf_mux_scbd_1793_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1793_up", this);
    pf_vf_mux_scbd_1794_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1794_up", this);
    pf_vf_mux_scbd_1795_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1795_up", this);
    pf_vf_mux_scbd_1796_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1796_up", this);
    pf_vf_mux_scbd_1797_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1797_up", this);
    pf_vf_mux_scbd_1798_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1798_up", this);
    pf_vf_mux_scbd_1799_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1799_up", this);
    pf_vf_mux_scbd_1800_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1800_up", this);
    pf_vf_mux_scbd_1801_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1801_up", this);
    pf_vf_mux_scbd_1802_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1802_up", this);
    pf_vf_mux_scbd_1803_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1803_up", this);
    pf_vf_mux_scbd_1804_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1804_up", this);
    pf_vf_mux_scbd_1805_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1805_up", this);
    pf_vf_mux_scbd_1806_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1806_up", this);
    pf_vf_mux_scbd_1807_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1807_up", this);
    pf_vf_mux_scbd_1808_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1808_up", this);
    pf_vf_mux_scbd_1809_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1809_up", this);
    pf_vf_mux_scbd_1810_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1810_up", this);
    pf_vf_mux_scbd_1811_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1811_up", this);
    pf_vf_mux_scbd_1812_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1812_up", this);
    pf_vf_mux_scbd_1813_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1813_up", this);
    pf_vf_mux_scbd_1814_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1814_up", this);
    pf_vf_mux_scbd_1815_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1815_up", this);
    pf_vf_mux_scbd_1816_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1816_up", this);
    pf_vf_mux_scbd_1817_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1817_up", this);
    pf_vf_mux_scbd_1818_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1818_up", this);
    pf_vf_mux_scbd_1819_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1819_up", this);
    pf_vf_mux_scbd_1820_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1820_up", this);
    pf_vf_mux_scbd_1821_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1821_up", this);
    pf_vf_mux_scbd_1822_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1822_up", this);
    pf_vf_mux_scbd_1823_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1823_up", this);
    pf_vf_mux_scbd_1824_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1824_up", this);
    pf_vf_mux_scbd_1825_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1825_up", this);
    pf_vf_mux_scbd_1826_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1826_up", this);
    pf_vf_mux_scbd_1827_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1827_up", this);
    pf_vf_mux_scbd_1828_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1828_up", this);
    pf_vf_mux_scbd_1829_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1829_up", this);
    pf_vf_mux_scbd_1830_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1830_up", this);
    pf_vf_mux_scbd_1831_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1831_up", this);
    pf_vf_mux_scbd_1832_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1832_up", this);
    pf_vf_mux_scbd_1833_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1833_up", this);
    pf_vf_mux_scbd_1834_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1834_up", this);
    pf_vf_mux_scbd_1835_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1835_up", this);
    pf_vf_mux_scbd_1836_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1836_up", this);
    pf_vf_mux_scbd_1837_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1837_up", this);
    pf_vf_mux_scbd_1838_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1838_up", this);
    pf_vf_mux_scbd_1839_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1839_up", this);
    pf_vf_mux_scbd_1840_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1840_up", this);
    pf_vf_mux_scbd_1841_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1841_up", this);
    pf_vf_mux_scbd_1842_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1842_up", this);
    pf_vf_mux_scbd_1843_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1843_up", this);
    pf_vf_mux_scbd_1844_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1844_up", this);
    pf_vf_mux_scbd_1845_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1845_up", this);
    pf_vf_mux_scbd_1846_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1846_up", this);
    pf_vf_mux_scbd_1847_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1847_up", this);
    pf_vf_mux_scbd_1848_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1848_up", this);
    pf_vf_mux_scbd_1849_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1849_up", this);
    pf_vf_mux_scbd_1850_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1850_up", this);
    pf_vf_mux_scbd_1851_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1851_up", this);
    pf_vf_mux_scbd_1852_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1852_up", this);
    pf_vf_mux_scbd_1853_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1853_up", this);
    pf_vf_mux_scbd_1854_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1854_up", this);
    pf_vf_mux_scbd_1855_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1855_up", this);
    pf_vf_mux_scbd_1856_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1856_up", this);
    pf_vf_mux_scbd_1857_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1857_up", this);
    pf_vf_mux_scbd_1858_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1858_up", this);
    pf_vf_mux_scbd_1859_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1859_up", this);
    pf_vf_mux_scbd_1860_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1860_up", this);
    pf_vf_mux_scbd_1861_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1861_up", this);
    pf_vf_mux_scbd_1862_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1862_up", this);
    pf_vf_mux_scbd_1863_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1863_up", this);
    pf_vf_mux_scbd_1864_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1864_up", this);
    pf_vf_mux_scbd_1865_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1865_up", this);
    pf_vf_mux_scbd_1866_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1866_up", this);
    pf_vf_mux_scbd_1867_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1867_up", this);
    pf_vf_mux_scbd_1868_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1868_up", this);
    pf_vf_mux_scbd_1869_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1869_up", this);
    pf_vf_mux_scbd_1870_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1870_up", this);
    pf_vf_mux_scbd_1871_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1871_up", this);
    pf_vf_mux_scbd_1872_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1872_up", this);
    pf_vf_mux_scbd_1873_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1873_up", this);
    pf_vf_mux_scbd_1874_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1874_up", this);
    pf_vf_mux_scbd_1875_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1875_up", this);
    pf_vf_mux_scbd_1876_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1876_up", this);
    pf_vf_mux_scbd_1877_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1877_up", this);
    pf_vf_mux_scbd_1878_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1878_up", this);
    pf_vf_mux_scbd_1879_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1879_up", this);
    pf_vf_mux_scbd_1880_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1880_up", this);
    pf_vf_mux_scbd_1881_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1881_up", this);
    pf_vf_mux_scbd_1882_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1882_up", this);
    pf_vf_mux_scbd_1883_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1883_up", this);
    pf_vf_mux_scbd_1884_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1884_up", this);
    pf_vf_mux_scbd_1885_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1885_up", this);
    pf_vf_mux_scbd_1886_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1886_up", this);
    pf_vf_mux_scbd_1887_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1887_up", this);
    pf_vf_mux_scbd_1888_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1888_up", this);
    pf_vf_mux_scbd_1889_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1889_up", this);
    pf_vf_mux_scbd_1890_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1890_up", this);
    pf_vf_mux_scbd_1891_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1891_up", this);
    pf_vf_mux_scbd_1892_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1892_up", this);
    pf_vf_mux_scbd_1893_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1893_up", this);
    pf_vf_mux_scbd_1894_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1894_up", this);
    pf_vf_mux_scbd_1895_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1895_up", this);
    pf_vf_mux_scbd_1896_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1896_up", this);
    pf_vf_mux_scbd_1897_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1897_up", this);
    pf_vf_mux_scbd_1898_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1898_up", this);
    pf_vf_mux_scbd_1899_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1899_up", this);
    pf_vf_mux_scbd_1900_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1900_up", this);
    pf_vf_mux_scbd_1901_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1901_up", this);
    pf_vf_mux_scbd_1902_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1902_up", this);
    pf_vf_mux_scbd_1903_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1903_up", this);
    pf_vf_mux_scbd_1904_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1904_up", this);
    pf_vf_mux_scbd_1905_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1905_up", this);
    pf_vf_mux_scbd_1906_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1906_up", this);
    pf_vf_mux_scbd_1907_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1907_up", this);
    pf_vf_mux_scbd_1908_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1908_up", this);
    pf_vf_mux_scbd_1909_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1909_up", this);
    pf_vf_mux_scbd_1910_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1910_up", this);
    pf_vf_mux_scbd_1911_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1911_up", this);
    pf_vf_mux_scbd_1912_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1912_up", this);
    pf_vf_mux_scbd_1913_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1913_up", this);
    pf_vf_mux_scbd_1914_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1914_up", this);
    pf_vf_mux_scbd_1915_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1915_up", this);
    pf_vf_mux_scbd_1916_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1916_up", this);
    pf_vf_mux_scbd_1917_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1917_up", this);
    pf_vf_mux_scbd_1918_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1918_up", this);
    pf_vf_mux_scbd_1919_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1919_up", this);
    pf_vf_mux_scbd_1920_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1920_up", this);
    pf_vf_mux_scbd_1921_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1921_up", this);
    pf_vf_mux_scbd_1922_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1922_up", this);
    pf_vf_mux_scbd_1923_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1923_up", this);
    pf_vf_mux_scbd_1924_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1924_up", this);
    pf_vf_mux_scbd_1925_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1925_up", this);
    pf_vf_mux_scbd_1926_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1926_up", this);
    pf_vf_mux_scbd_1927_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1927_up", this);
    pf_vf_mux_scbd_1928_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1928_up", this);
    pf_vf_mux_scbd_1929_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1929_up", this);
    pf_vf_mux_scbd_1930_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1930_up", this);
    pf_vf_mux_scbd_1931_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1931_up", this);
    pf_vf_mux_scbd_1932_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1932_up", this);
    pf_vf_mux_scbd_1933_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1933_up", this);
    pf_vf_mux_scbd_1934_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1934_up", this);
    pf_vf_mux_scbd_1935_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1935_up", this);
    pf_vf_mux_scbd_1936_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1936_up", this);
    pf_vf_mux_scbd_1937_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1937_up", this);
    pf_vf_mux_scbd_1938_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1938_up", this);
    pf_vf_mux_scbd_1939_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1939_up", this);
    pf_vf_mux_scbd_1940_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1940_up", this);
    pf_vf_mux_scbd_1941_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1941_up", this);
    pf_vf_mux_scbd_1942_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1942_up", this);
    pf_vf_mux_scbd_1943_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1943_up", this);
    pf_vf_mux_scbd_1944_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1944_up", this);
    pf_vf_mux_scbd_1945_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1945_up", this);
    pf_vf_mux_scbd_1946_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1946_up", this);
    pf_vf_mux_scbd_1947_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1947_up", this);
    pf_vf_mux_scbd_1948_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1948_up", this);
    pf_vf_mux_scbd_1949_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1949_up", this);
    pf_vf_mux_scbd_1950_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1950_up", this);
    pf_vf_mux_scbd_1951_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1951_up", this);
    pf_vf_mux_scbd_1952_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1952_up", this);
    pf_vf_mux_scbd_1953_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1953_up", this);
    pf_vf_mux_scbd_1954_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1954_up", this);
    pf_vf_mux_scbd_1955_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1955_up", this);
    pf_vf_mux_scbd_1956_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1956_up", this);
    pf_vf_mux_scbd_1957_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1957_up", this);
    pf_vf_mux_scbd_1958_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1958_up", this);
    pf_vf_mux_scbd_1959_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1959_up", this);
    pf_vf_mux_scbd_1960_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1960_up", this);
    pf_vf_mux_scbd_1961_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1961_up", this);
    pf_vf_mux_scbd_1962_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1962_up", this);
    pf_vf_mux_scbd_1963_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1963_up", this);
    pf_vf_mux_scbd_1964_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1964_up", this);
    pf_vf_mux_scbd_1965_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1965_up", this);
    pf_vf_mux_scbd_1966_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1966_up", this);
    pf_vf_mux_scbd_1967_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1967_up", this);
    pf_vf_mux_scbd_1968_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1968_up", this);
    pf_vf_mux_scbd_1969_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1969_up", this);
    pf_vf_mux_scbd_1970_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1970_up", this);
    pf_vf_mux_scbd_1971_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1971_up", this);
    pf_vf_mux_scbd_1972_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1972_up", this);
    pf_vf_mux_scbd_1973_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1973_up", this);
    pf_vf_mux_scbd_1974_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1974_up", this);
    pf_vf_mux_scbd_1975_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1975_up", this);
    pf_vf_mux_scbd_1976_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1976_up", this);
    pf_vf_mux_scbd_1977_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1977_up", this);
    pf_vf_mux_scbd_1978_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1978_up", this);
    pf_vf_mux_scbd_1979_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1979_up", this);
    pf_vf_mux_scbd_1980_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1980_up", this);
    pf_vf_mux_scbd_1981_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1981_up", this);
    pf_vf_mux_scbd_1982_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1982_up", this);
    pf_vf_mux_scbd_1983_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1983_up", this);
    pf_vf_mux_scbd_1984_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1984_up", this);
    pf_vf_mux_scbd_1985_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1985_up", this);
    pf_vf_mux_scbd_1986_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1986_up", this);
    pf_vf_mux_scbd_1987_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1987_up", this);
    pf_vf_mux_scbd_1988_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1988_up", this);
    pf_vf_mux_scbd_1989_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1989_up", this);
    pf_vf_mux_scbd_1990_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1990_up", this);
    pf_vf_mux_scbd_1991_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1991_up", this);
    pf_vf_mux_scbd_1992_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1992_up", this);
    pf_vf_mux_scbd_1993_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1993_up", this);
    pf_vf_mux_scbd_1994_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1994_up", this);
    pf_vf_mux_scbd_1995_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1995_up", this);
    pf_vf_mux_scbd_1996_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1996_up", this);
    pf_vf_mux_scbd_1997_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1997_up", this);
    pf_vf_mux_scbd_1998_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1998_up", this);
    pf_vf_mux_scbd_1999_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_1999_up", this);
    pf_vf_mux_scbd_2000_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2000_up", this);
    pf_vf_mux_scbd_2001_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2001_up", this);
    pf_vf_mux_scbd_2002_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2002_up", this);
    pf_vf_mux_scbd_2003_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2003_up", this);
    pf_vf_mux_scbd_2004_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2004_up", this);
    pf_vf_mux_scbd_2005_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2005_up", this);
    pf_vf_mux_scbd_2006_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2006_up", this);
    pf_vf_mux_scbd_2007_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2007_up", this);
    pf_vf_mux_scbd_2008_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2008_up", this);
    pf_vf_mux_scbd_2009_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2009_up", this);
    pf_vf_mux_scbd_2010_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2010_up", this);
    pf_vf_mux_scbd_2011_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2011_up", this);
    pf_vf_mux_scbd_2012_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2012_up", this);
    pf_vf_mux_scbd_2013_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2013_up", this);
    pf_vf_mux_scbd_2014_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2014_up", this);
    pf_vf_mux_scbd_2015_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2015_up", this);
    pf_vf_mux_scbd_2016_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2016_up", this);
    pf_vf_mux_scbd_2017_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2017_up", this);
    pf_vf_mux_scbd_2018_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2018_up", this);
    pf_vf_mux_scbd_2019_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2019_up", this);
    pf_vf_mux_scbd_2020_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2020_up", this);
    pf_vf_mux_scbd_2021_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2021_up", this);
    pf_vf_mux_scbd_2022_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2022_up", this);
    pf_vf_mux_scbd_2023_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2023_up", this);
    pf_vf_mux_scbd_2024_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2024_up", this);
    pf_vf_mux_scbd_2025_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2025_up", this);
    pf_vf_mux_scbd_2026_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2026_up", this);
    pf_vf_mux_scbd_2027_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2027_up", this);
    pf_vf_mux_scbd_2028_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2028_up", this);
    pf_vf_mux_scbd_2029_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2029_up", this);
    pf_vf_mux_scbd_2030_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2030_up", this);
    pf_vf_mux_scbd_2031_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2031_up", this);
    pf_vf_mux_scbd_2032_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2032_up", this);
    pf_vf_mux_scbd_2033_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2033_up", this);
    pf_vf_mux_scbd_2034_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2034_up", this);
    pf_vf_mux_scbd_2035_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2035_up", this);
    pf_vf_mux_scbd_2036_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2036_up", this);
    pf_vf_mux_scbd_2037_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2037_up", this);
    pf_vf_mux_scbd_2038_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2038_up", this);
    pf_vf_mux_scbd_2039_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2039_up", this);
    pf_vf_mux_scbd_2040_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2040_up", this);
    pf_vf_mux_scbd_2041_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2041_up", this);
    pf_vf_mux_scbd_2042_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2042_up", this);
    pf_vf_mux_scbd_2043_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2043_up", this);
    pf_vf_mux_scbd_2044_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2044_up", this);
    pf_vf_mux_scbd_2045_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2045_up", this);
    pf_vf_mux_scbd_2046_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2046_up", this);
    pf_vf_mux_scbd_2047_up = pf_vf_mux_scoreboard::type_id::create("pf_vf_mux_scbd_2047_up", this);


    `endif


    /** Construct the virtual sequencer */
    sequencer = pf_vf_mux_virtual_sequencer::type_id::create("sequencer", this);

    `uvm_info("build_phase", "Exiting...", UVM_LOW)
  endfunction

  // Connect master analysis ports to scoreboard
  function void connect_phase(uvm_phase phase);
    `uvm_info("connect_phase", "Entered...",UVM_LOW)

    `monitor_scoreboard_connection(0);
    `monitor_scoreboard_connection(1);
    `monitor_scoreboard_connection(2);
    `monitor_scoreboard_connection(3);
    `monitor_scoreboard_connection(4);
    `monitor_scoreboard_connection(5);
    `monitor_scoreboard_connection(6);
    `monitor_scoreboard_connection(7);
    `monitor_scoreboard_connection(8);
    `monitor_scoreboard_connection(9);
    `monitor_scoreboard_connection(10);
    `monitor_scoreboard_connection(11);
    `monitor_scoreboard_connection(12);
    `monitor_scoreboard_connection(13);
    `monitor_scoreboard_connection(14);
    `monitor_scoreboard_connection(15);
    `monitor_scoreboard_upstream_connection(0);
    `monitor_scoreboard_upstream_connection(1);
    `monitor_scoreboard_upstream_connection(2);
    `monitor_scoreboard_upstream_connection(3);
    `monitor_scoreboard_upstream_connection(4);
    `monitor_scoreboard_upstream_connection(5);
    `monitor_scoreboard_upstream_connection(6);
    `monitor_scoreboard_upstream_connection(7);
    `monitor_scoreboard_upstream_connection(8);
    `monitor_scoreboard_upstream_connection(9);
    `monitor_scoreboard_upstream_connection(10);
    `monitor_scoreboard_upstream_connection(11);
    `monitor_scoreboard_upstream_connection(12);
    `monitor_scoreboard_upstream_connection(13);
    `monitor_scoreboard_upstream_connection(14);
    `monitor_scoreboard_upstream_connection(15);

    `ifdef TB_CONFIG_2
    `monitor_scoreboard_connection_N(0,16);
    `monitor_scoreboard_connection_N(1,17);
    `monitor_scoreboard_connection_N(2,18);
    `monitor_scoreboard_connection_N(3,19);
    `monitor_scoreboard_connection_N(4,20);
    `monitor_scoreboard_connection_N(5,21);
    `monitor_scoreboard_connection_N(6,22);
    `monitor_scoreboard_connection_N(7,23);
    `monitor_scoreboard_upstream_connection_N(0,16);
    `monitor_scoreboard_upstream_connection_N(1,17);
    `monitor_scoreboard_upstream_connection_N(2,18);
    `monitor_scoreboard_upstream_connection_N(3,19);
    `monitor_scoreboard_upstream_connection_N(4,20);
    `monitor_scoreboard_upstream_connection_N(5,21);
    `monitor_scoreboard_upstream_connection_N(6,22);
    `monitor_scoreboard_upstream_connection_N(7,23);
    `elsif TB_CONFIG_3
    `monitor_scoreboard_connection_N(0,16);
    `monitor_scoreboard_connection_N(1,17);
    `monitor_scoreboard_connection_N(2,18);
    `monitor_scoreboard_connection_N(3,19);
    `monitor_scoreboard_connection_N(4,20);
    `monitor_scoreboard_connection_N(5,21);
    `monitor_scoreboard_connection_N(6,22);
    `monitor_scoreboard_connection_N(7,23);
    `monitor_scoreboard_connection_N(8,24);
    `monitor_scoreboard_connection_N(9,25);
    `monitor_scoreboard_connection_N(10,26);
    `monitor_scoreboard_connection_N(11,27);
    `monitor_scoreboard_connection_N(12,28);
    `monitor_scoreboard_connection_N(13,29);
    `monitor_scoreboard_connection_N(14,30);
    `monitor_scoreboard_connection_N(15,31);
    `monitor_scoreboard_upstream_connection_N(0,16);
    `monitor_scoreboard_upstream_connection_N(1,17);
    `monitor_scoreboard_upstream_connection_N(2,18);
    `monitor_scoreboard_upstream_connection_N(3,19);
    `monitor_scoreboard_upstream_connection_N(4,20);
    `monitor_scoreboard_upstream_connection_N(5,21);
    `monitor_scoreboard_upstream_connection_N(6,22);
    `monitor_scoreboard_upstream_connection_N(7,23);
    `monitor_scoreboard_upstream_connection_N(8,24);
    `monitor_scoreboard_upstream_connection_N(9,25);
    `monitor_scoreboard_upstream_connection_N(10,26);
    `monitor_scoreboard_upstream_connection_N(11,27);
    `monitor_scoreboard_upstream_connection_N(12,28);
    `monitor_scoreboard_upstream_connection_N(13,29);
    `monitor_scoreboard_upstream_connection_N(14,30);
    `monitor_scoreboard_upstream_connection_N(15,31);
    `elsif TB_CONFIG_4
    `monitor_scoreboard_connection(16);
    `monitor_scoreboard_connection(17);
    `monitor_scoreboard_connection(18);
    `monitor_scoreboard_connection(19);
    `monitor_scoreboard_connection(20);
    `monitor_scoreboard_connection(21);
    `monitor_scoreboard_connection(22);
    `monitor_scoreboard_connection(23);
    `monitor_scoreboard_connection(24);
    `monitor_scoreboard_connection(25);
    `monitor_scoreboard_connection(26);
    `monitor_scoreboard_connection(27);
    `monitor_scoreboard_connection(28);
    `monitor_scoreboard_connection(29);
    `monitor_scoreboard_connection(30);
    `monitor_scoreboard_connection(31);
    `monitor_scoreboard_connection(32);
    `monitor_scoreboard_connection(33);
    `monitor_scoreboard_connection(34);
    `monitor_scoreboard_connection(35);
    `monitor_scoreboard_connection(36);
    `monitor_scoreboard_connection(37);
    `monitor_scoreboard_connection(38);
    `monitor_scoreboard_connection(39);
    `monitor_scoreboard_connection(40);
    `monitor_scoreboard_connection(41);
    `monitor_scoreboard_connection(42);
    `monitor_scoreboard_connection(43);
    `monitor_scoreboard_connection(44);
    `monitor_scoreboard_connection(45);
    `monitor_scoreboard_connection(46);
    `monitor_scoreboard_connection(47);
    `monitor_scoreboard_connection(48);
    `monitor_scoreboard_connection(49);
    `monitor_scoreboard_connection(50);
    `monitor_scoreboard_connection(51);
    `monitor_scoreboard_connection(52);
    `monitor_scoreboard_connection(53);
    `monitor_scoreboard_connection(54);
    `monitor_scoreboard_connection(55);
    `monitor_scoreboard_connection(56);
    `monitor_scoreboard_connection(57);
    `monitor_scoreboard_connection(58);
    `monitor_scoreboard_connection(59);
    `monitor_scoreboard_connection(60);
    `monitor_scoreboard_connection(61);
    `monitor_scoreboard_connection(62);
    `monitor_scoreboard_connection(63);
    `monitor_scoreboard_connection(64);
    `monitor_scoreboard_connection(65);
    `monitor_scoreboard_connection(66);
    `monitor_scoreboard_connection(67);
    `monitor_scoreboard_connection(68);
    `monitor_scoreboard_connection(69);
    `monitor_scoreboard_connection(70);
    `monitor_scoreboard_connection(71);
    `monitor_scoreboard_connection(72);
    `monitor_scoreboard_connection(73);
    `monitor_scoreboard_connection(74);
    `monitor_scoreboard_connection(75);
    `monitor_scoreboard_connection(76);
    `monitor_scoreboard_connection(77);
    `monitor_scoreboard_connection(78);
    `monitor_scoreboard_connection(79);
    `monitor_scoreboard_connection(80);
    `monitor_scoreboard_connection(81);
    `monitor_scoreboard_connection(82);
    `monitor_scoreboard_connection(83);
    `monitor_scoreboard_connection(84);
    `monitor_scoreboard_connection(85);
    `monitor_scoreboard_connection(86);
    `monitor_scoreboard_connection(87);
    `monitor_scoreboard_connection(88);
    `monitor_scoreboard_connection(89);
    `monitor_scoreboard_connection(90);
    `monitor_scoreboard_connection(91);
    `monitor_scoreboard_connection(92);
    `monitor_scoreboard_connection(93);
    `monitor_scoreboard_connection(94);
    `monitor_scoreboard_connection(95);
    `monitor_scoreboard_connection(96);
    `monitor_scoreboard_connection(97);
    `monitor_scoreboard_connection(98);
    `monitor_scoreboard_connection(99);
    `monitor_scoreboard_connection(100);
    `monitor_scoreboard_connection(101);
    `monitor_scoreboard_connection(102);
    `monitor_scoreboard_connection(103);
    `monitor_scoreboard_connection(104);
    `monitor_scoreboard_connection(105);
    `monitor_scoreboard_connection(106);
    `monitor_scoreboard_connection(107);
    `monitor_scoreboard_connection(108);
    `monitor_scoreboard_connection(109);
    `monitor_scoreboard_connection(110);
    `monitor_scoreboard_connection(111);
    `monitor_scoreboard_connection(112);
    `monitor_scoreboard_connection(113);
    `monitor_scoreboard_connection(114);
    `monitor_scoreboard_connection(115);
    `monitor_scoreboard_connection(116);
    `monitor_scoreboard_connection(117);
    `monitor_scoreboard_connection(118);
    `monitor_scoreboard_connection(119);
    `monitor_scoreboard_connection(120);
    `monitor_scoreboard_connection(121);
    `monitor_scoreboard_connection(122);
    `monitor_scoreboard_connection(123);
    `monitor_scoreboard_connection(124);
    `monitor_scoreboard_connection(125);
    `monitor_scoreboard_connection(126);
    `monitor_scoreboard_connection(127);
    `monitor_scoreboard_connection(128);
    `monitor_scoreboard_connection(129);
    `monitor_scoreboard_connection(130);
    `monitor_scoreboard_connection(131);
    `monitor_scoreboard_connection(132);
    `monitor_scoreboard_connection(133);
    `monitor_scoreboard_connection(134);
    `monitor_scoreboard_connection(135);
    `monitor_scoreboard_connection(136);
    `monitor_scoreboard_connection(137);
    `monitor_scoreboard_connection(138);
    `monitor_scoreboard_connection(139);
    `monitor_scoreboard_connection(140);
    `monitor_scoreboard_connection(141);
    `monitor_scoreboard_connection(142);
    `monitor_scoreboard_connection(143);
    `monitor_scoreboard_connection(144);
    `monitor_scoreboard_connection(145);
    `monitor_scoreboard_connection(146);
    `monitor_scoreboard_connection(147);
    `monitor_scoreboard_connection(148);
    `monitor_scoreboard_connection(149);
    `monitor_scoreboard_connection(150);
    `monitor_scoreboard_connection(151);
    `monitor_scoreboard_connection(152);
    `monitor_scoreboard_connection(153);
    `monitor_scoreboard_connection(154);
    `monitor_scoreboard_connection(155);
    `monitor_scoreboard_connection(156);
    `monitor_scoreboard_connection(157);
    `monitor_scoreboard_connection(158);
    `monitor_scoreboard_connection(159);
    `monitor_scoreboard_connection(160);
    `monitor_scoreboard_connection(161);
    `monitor_scoreboard_connection(162);
    `monitor_scoreboard_connection(163);
    `monitor_scoreboard_connection(164);
    `monitor_scoreboard_connection(165);
    `monitor_scoreboard_connection(166);
    `monitor_scoreboard_connection(167);
    `monitor_scoreboard_connection(168);
    `monitor_scoreboard_connection(169);
    `monitor_scoreboard_connection(170);
    `monitor_scoreboard_connection(171);
    `monitor_scoreboard_connection(172);
    `monitor_scoreboard_connection(173);
    `monitor_scoreboard_connection(174);
    `monitor_scoreboard_connection(175);
    `monitor_scoreboard_connection(176);
    `monitor_scoreboard_connection(177);
    `monitor_scoreboard_connection(178);
    `monitor_scoreboard_connection(179);
    `monitor_scoreboard_connection(180);
    `monitor_scoreboard_connection(181);
    `monitor_scoreboard_connection(182);
    `monitor_scoreboard_connection(183);
    `monitor_scoreboard_connection(184);
    `monitor_scoreboard_connection(185);
    `monitor_scoreboard_connection(186);
    `monitor_scoreboard_connection(187);
    `monitor_scoreboard_connection(188);
    `monitor_scoreboard_connection(189);
    `monitor_scoreboard_connection(190);
    `monitor_scoreboard_connection(191);
    `monitor_scoreboard_connection(192);
    `monitor_scoreboard_connection(193);
    `monitor_scoreboard_connection(194);
    `monitor_scoreboard_connection(195);
    `monitor_scoreboard_connection(196);
    `monitor_scoreboard_connection(197);
    `monitor_scoreboard_connection(198);
    `monitor_scoreboard_connection(199);
    `monitor_scoreboard_connection(200);
    `monitor_scoreboard_connection(201);
    `monitor_scoreboard_connection(202);
    `monitor_scoreboard_connection(203);
    `monitor_scoreboard_connection(204);
    `monitor_scoreboard_connection(205);
    `monitor_scoreboard_connection(206);
    `monitor_scoreboard_connection(207);
    `monitor_scoreboard_connection(208);
    `monitor_scoreboard_connection(209);
    `monitor_scoreboard_connection(210);
    `monitor_scoreboard_connection(211);
    `monitor_scoreboard_connection(212);
    `monitor_scoreboard_connection(213);
    `monitor_scoreboard_connection(214);
    `monitor_scoreboard_connection(215);
    `monitor_scoreboard_connection(216);
    `monitor_scoreboard_connection(217);
    `monitor_scoreboard_connection(218);
    `monitor_scoreboard_connection(219);
    `monitor_scoreboard_connection(220);
    `monitor_scoreboard_connection(221);
    `monitor_scoreboard_connection(222);
    `monitor_scoreboard_connection(223);
    `monitor_scoreboard_connection(224);
    `monitor_scoreboard_connection(225);
    `monitor_scoreboard_connection(226);
    `monitor_scoreboard_connection(227);
    `monitor_scoreboard_connection(228);
    `monitor_scoreboard_connection(229);
    `monitor_scoreboard_connection(230);
    `monitor_scoreboard_connection(231);
    `monitor_scoreboard_connection(232);
    `monitor_scoreboard_connection(233);
    `monitor_scoreboard_connection(234);
    `monitor_scoreboard_connection(235);
    `monitor_scoreboard_connection(236);
    `monitor_scoreboard_connection(237);
    `monitor_scoreboard_connection(238);
    `monitor_scoreboard_connection(239);
    `monitor_scoreboard_connection(240);
    `monitor_scoreboard_connection(241);
    `monitor_scoreboard_connection(242);
    `monitor_scoreboard_connection(243);
    `monitor_scoreboard_connection(244);
    `monitor_scoreboard_connection(245);
    `monitor_scoreboard_connection(246);
    `monitor_scoreboard_connection(247);
    `monitor_scoreboard_connection(248);
    `monitor_scoreboard_connection(249);
    `monitor_scoreboard_connection(250);
    `monitor_scoreboard_connection(251);
    `monitor_scoreboard_connection(252);
    `monitor_scoreboard_connection(253);
    `monitor_scoreboard_connection(254);
    `monitor_scoreboard_connection(255);
    `monitor_scoreboard_connection(256);
    `monitor_scoreboard_connection(257);
    `monitor_scoreboard_connection(258);
    `monitor_scoreboard_connection(259);
    `monitor_scoreboard_connection(260);
    `monitor_scoreboard_connection(261);
    `monitor_scoreboard_connection(262);
    `monitor_scoreboard_connection(263);
    `monitor_scoreboard_connection(264);
    `monitor_scoreboard_connection(265);
    `monitor_scoreboard_connection(266);
    `monitor_scoreboard_connection(267);
    `monitor_scoreboard_connection(268);
    `monitor_scoreboard_connection(269);
    `monitor_scoreboard_connection(270);
    `monitor_scoreboard_connection(271);
    `monitor_scoreboard_connection(272);
    `monitor_scoreboard_connection(273);
    `monitor_scoreboard_connection(274);
    `monitor_scoreboard_connection(275);
    `monitor_scoreboard_connection(276);
    `monitor_scoreboard_connection(277);
    `monitor_scoreboard_connection(278);
    `monitor_scoreboard_connection(279);
    `monitor_scoreboard_connection(280);
    `monitor_scoreboard_connection(281);
    `monitor_scoreboard_connection(282);
    `monitor_scoreboard_connection(283);
    `monitor_scoreboard_connection(284);
    `monitor_scoreboard_connection(285);
    `monitor_scoreboard_connection(286);
    `monitor_scoreboard_connection(287);
    `monitor_scoreboard_connection(288);
    `monitor_scoreboard_connection(289);
    `monitor_scoreboard_connection(290);
    `monitor_scoreboard_connection(291);
    `monitor_scoreboard_connection(292);
    `monitor_scoreboard_connection(293);
    `monitor_scoreboard_connection(294);
    `monitor_scoreboard_connection(295);
    `monitor_scoreboard_connection(296);
    `monitor_scoreboard_connection(297);
    `monitor_scoreboard_connection(298);
    `monitor_scoreboard_connection(299);
    `monitor_scoreboard_connection(300);
    `monitor_scoreboard_connection(301);
    `monitor_scoreboard_connection(302);
    `monitor_scoreboard_connection(303);
    `monitor_scoreboard_connection(304);
    `monitor_scoreboard_connection(305);
    `monitor_scoreboard_connection(306);
    `monitor_scoreboard_connection(307);
    `monitor_scoreboard_connection(308);
    `monitor_scoreboard_connection(309);
    `monitor_scoreboard_connection(310);
    `monitor_scoreboard_connection(311);
    `monitor_scoreboard_connection(312);
    `monitor_scoreboard_connection(313);
    `monitor_scoreboard_connection(314);
    `monitor_scoreboard_connection(315);
    `monitor_scoreboard_connection(316);
    `monitor_scoreboard_connection(317);
    `monitor_scoreboard_connection(318);
    `monitor_scoreboard_connection(319);
    `monitor_scoreboard_connection(320);
    `monitor_scoreboard_connection(321);
    `monitor_scoreboard_connection(322);
    `monitor_scoreboard_connection(323);
    `monitor_scoreboard_connection(324);
    `monitor_scoreboard_connection(325);
    `monitor_scoreboard_connection(326);
    `monitor_scoreboard_connection(327);
    `monitor_scoreboard_connection(328);
    `monitor_scoreboard_connection(329);
    `monitor_scoreboard_connection(330);
    `monitor_scoreboard_connection(331);
    `monitor_scoreboard_connection(332);
    `monitor_scoreboard_connection(333);
    `monitor_scoreboard_connection(334);
    `monitor_scoreboard_connection(335);
    `monitor_scoreboard_connection(336);
    `monitor_scoreboard_connection(337);
    `monitor_scoreboard_connection(338);
    `monitor_scoreboard_connection(339);
    `monitor_scoreboard_connection(340);
    `monitor_scoreboard_connection(341);
    `monitor_scoreboard_connection(342);
    `monitor_scoreboard_connection(343);
    `monitor_scoreboard_connection(344);
    `monitor_scoreboard_connection(345);
    `monitor_scoreboard_connection(346);
    `monitor_scoreboard_connection(347);
    `monitor_scoreboard_connection(348);
    `monitor_scoreboard_connection(349);
    `monitor_scoreboard_connection(350);
    `monitor_scoreboard_connection(351);
    `monitor_scoreboard_connection(352);
    `monitor_scoreboard_connection(353);
    `monitor_scoreboard_connection(354);
    `monitor_scoreboard_connection(355);
    `monitor_scoreboard_connection(356);
    `monitor_scoreboard_connection(357);
    `monitor_scoreboard_connection(358);
    `monitor_scoreboard_connection(359);
    `monitor_scoreboard_connection(360);
    `monitor_scoreboard_connection(361);
    `monitor_scoreboard_connection(362);
    `monitor_scoreboard_connection(363);
    `monitor_scoreboard_connection(364);
    `monitor_scoreboard_connection(365);
    `monitor_scoreboard_connection(366);
    `monitor_scoreboard_connection(367);
    `monitor_scoreboard_connection(368);
    `monitor_scoreboard_connection(369);
    `monitor_scoreboard_connection(370);
    `monitor_scoreboard_connection(371);
    `monitor_scoreboard_connection(372);
    `monitor_scoreboard_connection(373);
    `monitor_scoreboard_connection(374);
    `monitor_scoreboard_connection(375);
    `monitor_scoreboard_connection(376);
    `monitor_scoreboard_connection(377);
    `monitor_scoreboard_connection(378);
    `monitor_scoreboard_connection(379);
    `monitor_scoreboard_connection(380);
    `monitor_scoreboard_connection(381);
    `monitor_scoreboard_connection(382);
    `monitor_scoreboard_connection(383);
    `monitor_scoreboard_connection(384);
    `monitor_scoreboard_connection(385);
    `monitor_scoreboard_connection(386);
    `monitor_scoreboard_connection(387);
    `monitor_scoreboard_connection(388);
    `monitor_scoreboard_connection(389);
    `monitor_scoreboard_connection(390);
    `monitor_scoreboard_connection(391);
    `monitor_scoreboard_connection(392);
    `monitor_scoreboard_connection(393);
    `monitor_scoreboard_connection(394);
    `monitor_scoreboard_connection(395);
    `monitor_scoreboard_connection(396);
    `monitor_scoreboard_connection(397);
    `monitor_scoreboard_connection(398);
    `monitor_scoreboard_connection(399);
    `monitor_scoreboard_connection(400);
    `monitor_scoreboard_connection(401);
    `monitor_scoreboard_connection(402);
    `monitor_scoreboard_connection(403);
    `monitor_scoreboard_connection(404);
    `monitor_scoreboard_connection(405);
    `monitor_scoreboard_connection(406);
    `monitor_scoreboard_connection(407);
    `monitor_scoreboard_connection(408);
    `monitor_scoreboard_connection(409);
    `monitor_scoreboard_connection(410);
    `monitor_scoreboard_connection(411);
    `monitor_scoreboard_connection(412);
    `monitor_scoreboard_connection(413);
    `monitor_scoreboard_connection(414);
    `monitor_scoreboard_connection(415);
    `monitor_scoreboard_connection(416);
    `monitor_scoreboard_connection(417);
    `monitor_scoreboard_connection(418);
    `monitor_scoreboard_connection(419);
    `monitor_scoreboard_connection(420);
    `monitor_scoreboard_connection(421);
    `monitor_scoreboard_connection(422);
    `monitor_scoreboard_connection(423);
    `monitor_scoreboard_connection(424);
    `monitor_scoreboard_connection(425);
    `monitor_scoreboard_connection(426);
    `monitor_scoreboard_connection(427);
    `monitor_scoreboard_connection(428);
    `monitor_scoreboard_connection(429);
    `monitor_scoreboard_connection(430);
    `monitor_scoreboard_connection(431);
    `monitor_scoreboard_connection(432);
    `monitor_scoreboard_connection(433);
    `monitor_scoreboard_connection(434);
    `monitor_scoreboard_connection(435);
    `monitor_scoreboard_connection(436);
    `monitor_scoreboard_connection(437);
    `monitor_scoreboard_connection(438);
    `monitor_scoreboard_connection(439);
    `monitor_scoreboard_connection(440);
    `monitor_scoreboard_connection(441);
    `monitor_scoreboard_connection(442);
    `monitor_scoreboard_connection(443);
    `monitor_scoreboard_connection(444);
    `monitor_scoreboard_connection(445);
    `monitor_scoreboard_connection(446);
    `monitor_scoreboard_connection(447);
    `monitor_scoreboard_connection(448);
    `monitor_scoreboard_connection(449);
    `monitor_scoreboard_connection_TB4(0,450,0);
    `monitor_scoreboard_connection_TB4(0,451,1);
    `monitor_scoreboard_connection_TB4(0,452,2);
    `monitor_scoreboard_connection_TB4(0,453,3);
    `monitor_scoreboard_connection_TB4(0,454,4);
    `monitor_scoreboard_connection_TB4(0,455,5);
    `monitor_scoreboard_connection_TB4(0,456,6);
    `monitor_scoreboard_connection_TB4(0,457,7);
    `monitor_scoreboard_connection_TB4(0,458,8);
    `monitor_scoreboard_connection_TB4(0,459,9);
    `monitor_scoreboard_connection_TB4(0,460,10);
    `monitor_scoreboard_connection_TB4(0,461,11);
    `monitor_scoreboard_connection_TB4(0,462,12);
    `monitor_scoreboard_connection_TB4(0,463,13);
    `monitor_scoreboard_connection_TB4(0,464,14);
    `monitor_scoreboard_connection_TB4(0,465,15);
    `monitor_scoreboard_connection_TB4(0,466,16);
    `monitor_scoreboard_connection_TB4(0,467,17);
    `monitor_scoreboard_connection_TB4(0,468,18);
    `monitor_scoreboard_connection_TB4(0,469,19);
    `monitor_scoreboard_connection_TB4(0,470,20);
    `monitor_scoreboard_connection_TB4(0,471,21);
    `monitor_scoreboard_connection_TB4(0,472,22);
    `monitor_scoreboard_connection_TB4(0,473,23);
    `monitor_scoreboard_connection_TB4(0,474,24);
    `monitor_scoreboard_connection_TB4(0,475,25);
    `monitor_scoreboard_connection_TB4(0,476,26);
    `monitor_scoreboard_connection_TB4(0,477,27);
    `monitor_scoreboard_connection_TB4(0,478,28);
    `monitor_scoreboard_connection_TB4(0,479,29);
    `monitor_scoreboard_connection_TB4(0,480,30);
    `monitor_scoreboard_connection_TB4(0,481,31);
    `monitor_scoreboard_connection_TB4(0,482,32);
    `monitor_scoreboard_connection_TB4(0,483,33);
    `monitor_scoreboard_connection_TB4(0,484,34);
    `monitor_scoreboard_connection_TB4(0,485,35);
    `monitor_scoreboard_connection_TB4(0,486,36);
    `monitor_scoreboard_connection_TB4(0,487,37);
    `monitor_scoreboard_connection_TB4(0,488,38);
    `monitor_scoreboard_connection_TB4(0,489,39);
    `monitor_scoreboard_connection_TB4(0,490,40);
    `monitor_scoreboard_connection_TB4(0,491,41);
    `monitor_scoreboard_connection_TB4(0,492,42);
    `monitor_scoreboard_connection_TB4(0,493,43);
    `monitor_scoreboard_connection_TB4(0,494,44);
    `monitor_scoreboard_connection_TB4(0,495,45);
    `monitor_scoreboard_connection_TB4(0,496,46);
    `monitor_scoreboard_connection_TB4(0,497,47);
    `monitor_scoreboard_connection_TB4(0,498,48);
    `monitor_scoreboard_connection_TB4(0,499,49);
    `monitor_scoreboard_connection_TB4(0,500,50);
    `monitor_scoreboard_connection_TB4(0,501,51);
    `monitor_scoreboard_connection_TB4(0,502,52);
    `monitor_scoreboard_connection_TB4(0,503,53);
    `monitor_scoreboard_connection_TB4(0,504,54);
    `monitor_scoreboard_connection_TB4(0,505,55);
    `monitor_scoreboard_connection_TB4(0,506,56);
    `monitor_scoreboard_connection_TB4(0,507,57);
    `monitor_scoreboard_connection_TB4(0,508,58);
    `monitor_scoreboard_connection_TB4(0,509,59);
    `monitor_scoreboard_connection_TB4(0,510,60);
    `monitor_scoreboard_connection_TB4(0,511,61);
    `monitor_scoreboard_connection_TB4(0,512,62);
    `monitor_scoreboard_connection_TB4(0,513,63);
    `monitor_scoreboard_connection_TB4(0,514,64);
    `monitor_scoreboard_connection_TB4(0,515,65);
    `monitor_scoreboard_connection_TB4(0,516,66);
    `monitor_scoreboard_connection_TB4(0,517,67);
    `monitor_scoreboard_connection_TB4(0,518,68);
    `monitor_scoreboard_connection_TB4(0,519,69);
    `monitor_scoreboard_connection_TB4(0,520,70);
    `monitor_scoreboard_connection_TB4(0,521,71);
    `monitor_scoreboard_connection_TB4(0,522,72);
    `monitor_scoreboard_connection_TB4(0,523,73);
    `monitor_scoreboard_connection_TB4(0,524,74);
    `monitor_scoreboard_connection_TB4(0,525,75);
    `monitor_scoreboard_connection_TB4(0,526,76);
    `monitor_scoreboard_connection_TB4(0,527,77);
    `monitor_scoreboard_connection_TB4(0,528,78);
    `monitor_scoreboard_connection_TB4(0,529,79);
    `monitor_scoreboard_connection_TB4(0,530,80);
    `monitor_scoreboard_connection_TB4(0,531,81);
    `monitor_scoreboard_connection_TB4(0,532,82);
    `monitor_scoreboard_connection_TB4(0,533,83);
    `monitor_scoreboard_connection_TB4(0,534,84);
    `monitor_scoreboard_connection_TB4(0,535,85);
    `monitor_scoreboard_connection_TB4(0,536,86);
    `monitor_scoreboard_connection_TB4(0,537,87);
    `monitor_scoreboard_connection_TB4(0,538,88);
    `monitor_scoreboard_connection_TB4(0,539,89);
    `monitor_scoreboard_connection_TB4(0,540,90);
    `monitor_scoreboard_connection_TB4(0,541,91);
    `monitor_scoreboard_connection_TB4(0,542,92);
    `monitor_scoreboard_connection_TB4(0,543,93);
    `monitor_scoreboard_connection_TB4(0,544,94);
    `monitor_scoreboard_connection_TB4(0,545,95);
    `monitor_scoreboard_connection_TB4(0,546,96);
    `monitor_scoreboard_connection_TB4(0,547,97);
    `monitor_scoreboard_connection_TB4(0,548,98);
    `monitor_scoreboard_connection_TB4(0,549,99);
    `monitor_scoreboard_connection_TB4(0,550,100);
    `monitor_scoreboard_connection_TB4(0,551,101);
    `monitor_scoreboard_connection_TB4(0,552,102);
    `monitor_scoreboard_connection_TB4(0,553,103);
    `monitor_scoreboard_connection_TB4(0,554,104);
    `monitor_scoreboard_connection_TB4(0,555,105);
    `monitor_scoreboard_connection_TB4(0,556,106);
    `monitor_scoreboard_connection_TB4(0,557,107);
    `monitor_scoreboard_connection_TB4(0,558,108);
    `monitor_scoreboard_connection_TB4(0,559,109);
    `monitor_scoreboard_connection_TB4(0,560,110);
    `monitor_scoreboard_connection_TB4(0,561,111);
    `monitor_scoreboard_connection_TB4(0,562,112);
    `monitor_scoreboard_connection_TB4(0,563,113);
    `monitor_scoreboard_connection_TB4(0,564,114);
    `monitor_scoreboard_connection_TB4(0,565,115);
    `monitor_scoreboard_connection_TB4(0,566,116);
    `monitor_scoreboard_connection_TB4(0,567,117);
    `monitor_scoreboard_connection_TB4(0,568,118);
    `monitor_scoreboard_connection_TB4(0,569,119);
    `monitor_scoreboard_connection_TB4(0,570,120);
    `monitor_scoreboard_connection_TB4(0,571,121);
    `monitor_scoreboard_connection_TB4(0,572,122);
    `monitor_scoreboard_connection_TB4(0,573,123);
    `monitor_scoreboard_connection_TB4(0,574,124);
    `monitor_scoreboard_connection_TB4(0,575,125);
    `monitor_scoreboard_connection_TB4(0,576,126);
    `monitor_scoreboard_connection_TB4(0,577,127);
    `monitor_scoreboard_connection_TB4(0,578,128);
    `monitor_scoreboard_connection_TB4(0,579,129);
    `monitor_scoreboard_connection_TB4(0,580,130);
    `monitor_scoreboard_connection_TB4(0,581,131);
    `monitor_scoreboard_connection_TB4(0,582,132);
    `monitor_scoreboard_connection_TB4(0,583,133);
    `monitor_scoreboard_connection_TB4(0,584,134);
    `monitor_scoreboard_connection_TB4(0,585,135);
    `monitor_scoreboard_connection_TB4(0,586,136);
    `monitor_scoreboard_connection_TB4(0,587,137);
    `monitor_scoreboard_connection_TB4(0,588,138);
    `monitor_scoreboard_connection_TB4(0,589,139);
    `monitor_scoreboard_connection_TB4(0,590,140);
    `monitor_scoreboard_connection_TB4(0,591,141);
    `monitor_scoreboard_connection_TB4(0,592,142);
    `monitor_scoreboard_connection_TB4(0,593,143);
    `monitor_scoreboard_connection_TB4(0,594,144);
    `monitor_scoreboard_connection_TB4(0,595,145);
    `monitor_scoreboard_connection_TB4(0,596,146);
    `monitor_scoreboard_connection_TB4(0,597,147);
    `monitor_scoreboard_connection_TB4(0,598,148);
    `monitor_scoreboard_connection_TB4(0,599,149);
    `monitor_scoreboard_connection_TB4(0,600,150);
    `monitor_scoreboard_connection_TB4(0,601,151);
    `monitor_scoreboard_connection_TB4(0,602,152);
    `monitor_scoreboard_connection_TB4(0,603,153);
    `monitor_scoreboard_connection_TB4(0,604,154);
    `monitor_scoreboard_connection_TB4(0,605,155);
    `monitor_scoreboard_connection_TB4(0,606,156);
    `monitor_scoreboard_connection_TB4(0,607,157);
    `monitor_scoreboard_connection_TB4(0,608,158);
    `monitor_scoreboard_connection_TB4(0,609,159);
    `monitor_scoreboard_connection_TB4(0,610,160);
    `monitor_scoreboard_connection_TB4(0,611,161);
    `monitor_scoreboard_connection_TB4(0,612,162);
    `monitor_scoreboard_connection_TB4(0,613,163);
    `monitor_scoreboard_connection_TB4(0,614,164);
    `monitor_scoreboard_connection_TB4(0,615,165);
    `monitor_scoreboard_connection_TB4(0,616,166);
    `monitor_scoreboard_connection_TB4(0,617,167);
    `monitor_scoreboard_connection_TB4(0,618,168);
    `monitor_scoreboard_connection_TB4(0,619,169);
    `monitor_scoreboard_connection_TB4(0,620,170);
    `monitor_scoreboard_connection_TB4(0,621,171);
    `monitor_scoreboard_connection_TB4(0,622,172);
    `monitor_scoreboard_connection_TB4(0,623,173);
    `monitor_scoreboard_connection_TB4(0,624,174);
    `monitor_scoreboard_connection_TB4(0,625,175);
    `monitor_scoreboard_connection_TB4(0,626,176);
    `monitor_scoreboard_connection_TB4(0,627,177);
    `monitor_scoreboard_connection_TB4(0,628,178);
    `monitor_scoreboard_connection_TB4(0,629,179);
    `monitor_scoreboard_connection_TB4(0,630,180);
    `monitor_scoreboard_connection_TB4(0,631,181);
    `monitor_scoreboard_connection_TB4(0,632,182);
    `monitor_scoreboard_connection_TB4(0,633,183);
    `monitor_scoreboard_connection_TB4(0,634,184);
    `monitor_scoreboard_connection_TB4(0,635,185);
    `monitor_scoreboard_connection_TB4(0,636,186);
    `monitor_scoreboard_connection_TB4(0,637,187);
    `monitor_scoreboard_connection_TB4(0,638,188);
    `monitor_scoreboard_connection_TB4(0,639,189);
    `monitor_scoreboard_connection_TB4(0,640,190);
    `monitor_scoreboard_connection_TB4(0,641,191);
    `monitor_scoreboard_connection_TB4(0,642,192);
    `monitor_scoreboard_connection_TB4(0,643,193);
    `monitor_scoreboard_connection_TB4(0,644,194);
    `monitor_scoreboard_connection_TB4(0,645,195);
    `monitor_scoreboard_connection_TB4(0,646,196);
    `monitor_scoreboard_connection_TB4(0,647,197);
    `monitor_scoreboard_connection_TB4(0,648,198);
    `monitor_scoreboard_connection_TB4(0,649,199);
    `monitor_scoreboard_connection_TB4(0,650,200);
    `monitor_scoreboard_connection_TB4(0,651,201);
    `monitor_scoreboard_connection_TB4(0,652,202);
    `monitor_scoreboard_connection_TB4(0,653,203);
    `monitor_scoreboard_connection_TB4(0,654,204);
    `monitor_scoreboard_connection_TB4(0,655,205);
    `monitor_scoreboard_connection_TB4(0,656,206);
    `monitor_scoreboard_connection_TB4(0,657,207);
    `monitor_scoreboard_connection_TB4(0,658,208);
    `monitor_scoreboard_connection_TB4(0,659,209);
    `monitor_scoreboard_connection_TB4(0,660,210);
    `monitor_scoreboard_connection_TB4(0,661,211);
    `monitor_scoreboard_connection_TB4(0,662,212);
    `monitor_scoreboard_connection_TB4(0,663,213);
    `monitor_scoreboard_connection_TB4(0,664,214);
    `monitor_scoreboard_connection_TB4(0,665,215);
    `monitor_scoreboard_connection_TB4(0,666,216);
    `monitor_scoreboard_connection_TB4(0,667,217);
    `monitor_scoreboard_connection_TB4(0,668,218);
    `monitor_scoreboard_connection_TB4(0,669,219);
    `monitor_scoreboard_connection_TB4(0,670,220);
    `monitor_scoreboard_connection_TB4(0,671,221);
    `monitor_scoreboard_connection_TB4(0,672,222);
    `monitor_scoreboard_connection_TB4(0,673,223);
    `monitor_scoreboard_connection_TB4(0,674,224);
    `monitor_scoreboard_connection_TB4(0,675,225);
    `monitor_scoreboard_connection_TB4(0,676,226);
    `monitor_scoreboard_connection_TB4(0,677,227);
    `monitor_scoreboard_connection_TB4(0,678,228);
    `monitor_scoreboard_connection_TB4(0,679,229);
    `monitor_scoreboard_connection_TB4(0,680,230);
    `monitor_scoreboard_connection_TB4(0,681,231);
    `monitor_scoreboard_connection_TB4(0,682,232);
    `monitor_scoreboard_connection_TB4(0,683,233);
    `monitor_scoreboard_connection_TB4(0,684,234);
    `monitor_scoreboard_connection_TB4(0,685,235);
    `monitor_scoreboard_connection_TB4(0,686,236);
    `monitor_scoreboard_connection_TB4(0,687,237);
    `monitor_scoreboard_connection_TB4(0,688,238);
    `monitor_scoreboard_connection_TB4(0,689,239);
    `monitor_scoreboard_connection_TB4(0,690,240);
    `monitor_scoreboard_connection_TB4(0,691,241);
    `monitor_scoreboard_connection_TB4(0,692,242);
    `monitor_scoreboard_connection_TB4(0,693,243);
    `monitor_scoreboard_connection_TB4(0,694,244);
    `monitor_scoreboard_connection_TB4(0,695,245);
    `monitor_scoreboard_connection_TB4(0,696,246);
    `monitor_scoreboard_connection_TB4(0,697,247);
    `monitor_scoreboard_connection_TB4(0,698,248);
    `monitor_scoreboard_connection_TB4(0,699,249);
    `monitor_scoreboard_connection_TB4(0,700,250);
    `monitor_scoreboard_connection_TB4(0,701,251);
    `monitor_scoreboard_connection_TB4(0,702,252);
    `monitor_scoreboard_connection_TB4(0,703,253);
    `monitor_scoreboard_connection_TB4(0,704,254);
    `monitor_scoreboard_connection_TB4(0,705,255);
    `monitor_scoreboard_connection_TB4(0,706,256);
    `monitor_scoreboard_connection_TB4(0,707,257);
    `monitor_scoreboard_connection_TB4(0,708,258);
    `monitor_scoreboard_connection_TB4(0,709,259);
    `monitor_scoreboard_connection_TB4(0,710,260);
    `monitor_scoreboard_connection_TB4(0,711,261);
    `monitor_scoreboard_connection_TB4(0,712,262);
    `monitor_scoreboard_connection_TB4(0,713,263);
    `monitor_scoreboard_connection_TB4(0,714,264);
    `monitor_scoreboard_connection_TB4(0,715,265);
    `monitor_scoreboard_connection_TB4(0,716,266);
    `monitor_scoreboard_connection_TB4(0,717,267);
    `monitor_scoreboard_connection_TB4(0,718,268);
    `monitor_scoreboard_connection_TB4(0,719,269);
    `monitor_scoreboard_connection_TB4(0,720,270);
    `monitor_scoreboard_connection_TB4(0,721,271);
    `monitor_scoreboard_connection_TB4(0,722,272);
    `monitor_scoreboard_connection_TB4(0,723,273);
    `monitor_scoreboard_connection_TB4(0,724,274);
    `monitor_scoreboard_connection_TB4(0,725,275);
    `monitor_scoreboard_connection_TB4(0,726,276);
    `monitor_scoreboard_connection_TB4(0,727,277);
    `monitor_scoreboard_connection_TB4(0,728,278);
    `monitor_scoreboard_connection_TB4(0,729,279);
    `monitor_scoreboard_connection_TB4(0,730,280);
    `monitor_scoreboard_connection_TB4(0,731,281);
    `monitor_scoreboard_connection_TB4(0,732,282);
    `monitor_scoreboard_connection_TB4(0,733,283);
    `monitor_scoreboard_connection_TB4(0,734,284);
    `monitor_scoreboard_connection_TB4(0,735,285);
    `monitor_scoreboard_connection_TB4(0,736,286);
    `monitor_scoreboard_connection_TB4(0,737,287);
    `monitor_scoreboard_connection_TB4(0,738,288);
    `monitor_scoreboard_connection_TB4(0,739,289);
    `monitor_scoreboard_connection_TB4(0,740,290);
    `monitor_scoreboard_connection_TB4(0,741,291);
    `monitor_scoreboard_connection_TB4(0,742,292);
    `monitor_scoreboard_connection_TB4(0,743,293);
    `monitor_scoreboard_connection_TB4(0,744,294);
    `monitor_scoreboard_connection_TB4(0,745,295);
    `monitor_scoreboard_connection_TB4(0,746,296);
    `monitor_scoreboard_connection_TB4(0,747,297);
    `monitor_scoreboard_connection_TB4(0,748,298);
    `monitor_scoreboard_connection_TB4(0,749,299);
    `monitor_scoreboard_connection_TB4(0,750,300);
    `monitor_scoreboard_connection_TB4(0,751,301);
    `monitor_scoreboard_connection_TB4(0,752,302);
    `monitor_scoreboard_connection_TB4(0,753,303);
    `monitor_scoreboard_connection_TB4(0,754,304);
    `monitor_scoreboard_connection_TB4(0,755,305);
    `monitor_scoreboard_connection_TB4(0,756,306);
    `monitor_scoreboard_connection_TB4(0,757,307);
    `monitor_scoreboard_connection_TB4(0,758,308);
    `monitor_scoreboard_connection_TB4(0,759,309);
    `monitor_scoreboard_connection_TB4(0,760,310);
    `monitor_scoreboard_connection_TB4(0,761,311);
    `monitor_scoreboard_connection_TB4(0,762,312);
    `monitor_scoreboard_connection_TB4(0,763,313);
    `monitor_scoreboard_connection_TB4(0,764,314);
    `monitor_scoreboard_connection_TB4(0,765,315);
    `monitor_scoreboard_connection_TB4(0,766,316);
    `monitor_scoreboard_connection_TB4(0,767,317);
    `monitor_scoreboard_connection_TB4(0,768,318);
    `monitor_scoreboard_connection_TB4(0,769,319);
    `monitor_scoreboard_connection_TB4(0,770,320);
    `monitor_scoreboard_connection_TB4(0,771,321);
    `monitor_scoreboard_connection_TB4(0,772,322);
    `monitor_scoreboard_connection_TB4(0,773,323);
    `monitor_scoreboard_connection_TB4(0,774,324);
    `monitor_scoreboard_connection_TB4(0,775,325);
    `monitor_scoreboard_connection_TB4(0,776,326);
    `monitor_scoreboard_connection_TB4(0,777,327);
    `monitor_scoreboard_connection_TB4(0,778,328);
    `monitor_scoreboard_connection_TB4(0,779,329);
    `monitor_scoreboard_connection_TB4(0,780,330);
    `monitor_scoreboard_connection_TB4(0,781,331);
    `monitor_scoreboard_connection_TB4(0,782,332);
    `monitor_scoreboard_connection_TB4(0,783,333);
    `monitor_scoreboard_connection_TB4(0,784,334);
    `monitor_scoreboard_connection_TB4(0,785,335);
    `monitor_scoreboard_connection_TB4(0,786,336);
    `monitor_scoreboard_connection_TB4(0,787,337);
    `monitor_scoreboard_connection_TB4(0,788,338);
    `monitor_scoreboard_connection_TB4(0,789,339);
    `monitor_scoreboard_connection_TB4(0,790,340);
    `monitor_scoreboard_connection_TB4(0,791,341);
    `monitor_scoreboard_connection_TB4(0,792,342);
    `monitor_scoreboard_connection_TB4(0,793,343);
    `monitor_scoreboard_connection_TB4(0,794,344);
    `monitor_scoreboard_connection_TB4(0,795,345);
    `monitor_scoreboard_connection_TB4(0,796,346);
    `monitor_scoreboard_connection_TB4(0,797,347);
    `monitor_scoreboard_connection_TB4(0,798,348);
    `monitor_scoreboard_connection_TB4(0,799,349);
    `monitor_scoreboard_connection_TB4(0,800,350);
    `monitor_scoreboard_connection_TB4(0,801,351);
    `monitor_scoreboard_connection_TB4(0,802,352);
    `monitor_scoreboard_connection_TB4(0,803,353);
    `monitor_scoreboard_connection_TB4(0,804,354);
    `monitor_scoreboard_connection_TB4(0,805,355);
    `monitor_scoreboard_connection_TB4(0,806,356);
    `monitor_scoreboard_connection_TB4(0,807,357);
    `monitor_scoreboard_connection_TB4(0,808,358);
    `monitor_scoreboard_connection_TB4(0,809,359);
    `monitor_scoreboard_connection_TB4(0,810,360);
    `monitor_scoreboard_connection_TB4(0,811,361);
    `monitor_scoreboard_connection_TB4(0,812,362);
    `monitor_scoreboard_connection_TB4(0,813,363);
    `monitor_scoreboard_connection_TB4(0,814,364);
    `monitor_scoreboard_connection_TB4(0,815,365);
    `monitor_scoreboard_connection_TB4(0,816,366);
    `monitor_scoreboard_connection_TB4(0,817,367);
    `monitor_scoreboard_connection_TB4(0,818,368);
    `monitor_scoreboard_connection_TB4(0,819,369);
    `monitor_scoreboard_connection_TB4(0,820,370);
    `monitor_scoreboard_connection_TB4(0,821,371);
    `monitor_scoreboard_connection_TB4(0,822,372);
    `monitor_scoreboard_connection_TB4(0,823,373);
    `monitor_scoreboard_connection_TB4(0,824,374);
    `monitor_scoreboard_connection_TB4(0,825,375);
    `monitor_scoreboard_connection_TB4(0,826,376);
    `monitor_scoreboard_connection_TB4(0,827,377);
    `monitor_scoreboard_connection_TB4(0,828,378);
    `monitor_scoreboard_connection_TB4(0,829,379);
    `monitor_scoreboard_connection_TB4(0,830,380);
    `monitor_scoreboard_connection_TB4(0,831,381);
    `monitor_scoreboard_connection_TB4(0,832,382);
    `monitor_scoreboard_connection_TB4(0,833,383);
    `monitor_scoreboard_connection_TB4(0,834,384);
    `monitor_scoreboard_connection_TB4(0,835,385);
    `monitor_scoreboard_connection_TB4(0,836,386);
    `monitor_scoreboard_connection_TB4(0,837,387);
    `monitor_scoreboard_connection_TB4(0,838,388);
    `monitor_scoreboard_connection_TB4(0,839,389);
    `monitor_scoreboard_connection_TB4(0,840,390);
    `monitor_scoreboard_connection_TB4(0,841,391);
    `monitor_scoreboard_connection_TB4(0,842,392);
    `monitor_scoreboard_connection_TB4(0,843,393);
    `monitor_scoreboard_connection_TB4(0,844,394);
    `monitor_scoreboard_connection_TB4(0,845,395);
    `monitor_scoreboard_connection_TB4(0,846,396);
    `monitor_scoreboard_connection_TB4(0,847,397);
    `monitor_scoreboard_connection_TB4(0,848,398);
    `monitor_scoreboard_connection_TB4(0,849,399);
    `monitor_scoreboard_connection_TB4(0,850,400);
    `monitor_scoreboard_connection_TB4(0,851,401);
    `monitor_scoreboard_connection_TB4(0,852,402);
    `monitor_scoreboard_connection_TB4(0,853,403);
    `monitor_scoreboard_connection_TB4(0,854,404);
    `monitor_scoreboard_connection_TB4(0,855,405);
    `monitor_scoreboard_connection_TB4(0,856,406);
    `monitor_scoreboard_connection_TB4(0,857,407);
    `monitor_scoreboard_connection_TB4(0,858,408);
    `monitor_scoreboard_connection_TB4(0,859,409);
    `monitor_scoreboard_connection_TB4(0,860,410);
    `monitor_scoreboard_connection_TB4(0,861,411);
    `monitor_scoreboard_connection_TB4(0,862,412);
    `monitor_scoreboard_connection_TB4(0,863,413);
    `monitor_scoreboard_connection_TB4(0,864,414);
    `monitor_scoreboard_connection_TB4(0,865,415);
    `monitor_scoreboard_connection_TB4(0,866,416);
    `monitor_scoreboard_connection_TB4(0,867,417);
    `monitor_scoreboard_connection_TB4(0,868,418);
    `monitor_scoreboard_connection_TB4(0,869,419);
    `monitor_scoreboard_connection_TB4(0,870,420);
    `monitor_scoreboard_connection_TB4(0,871,421);
    `monitor_scoreboard_connection_TB4(0,872,422);
    `monitor_scoreboard_connection_TB4(0,873,423);
    `monitor_scoreboard_connection_TB4(0,874,424);
    `monitor_scoreboard_connection_TB4(0,875,425);
    `monitor_scoreboard_connection_TB4(0,876,426);
    `monitor_scoreboard_connection_TB4(0,877,427);
    `monitor_scoreboard_connection_TB4(0,878,428);
    `monitor_scoreboard_connection_TB4(0,879,429);
    `monitor_scoreboard_connection_TB4(0,880,430);
    `monitor_scoreboard_connection_TB4(0,881,431);
    `monitor_scoreboard_connection_TB4(0,882,432);
    `monitor_scoreboard_connection_TB4(0,883,433);
    `monitor_scoreboard_connection_TB4(0,884,434);
    `monitor_scoreboard_connection_TB4(0,885,435);
    `monitor_scoreboard_connection_TB4(0,886,436);
    `monitor_scoreboard_connection_TB4(0,887,437);
    `monitor_scoreboard_connection_TB4(0,888,438);
    `monitor_scoreboard_connection_TB4(0,889,439);
    `monitor_scoreboard_connection_TB4(0,890,440);
    `monitor_scoreboard_connection_TB4(0,891,441);
    `monitor_scoreboard_connection_TB4(0,892,442);
    `monitor_scoreboard_connection_TB4(0,893,443);
    `monitor_scoreboard_connection_TB4(0,894,444);
    `monitor_scoreboard_connection_TB4(0,895,445);
    `monitor_scoreboard_connection_TB4(0,896,446);
    `monitor_scoreboard_connection_TB4(0,897,447);
    `monitor_scoreboard_connection_TB4(0,898,448);
    `monitor_scoreboard_connection_TB4(0,899,449);
    `monitor_scoreboard_connection_TB4(1,900,0);
    `monitor_scoreboard_connection_TB4(1,901,1);
    `monitor_scoreboard_connection_TB4(1,902,2);
    `monitor_scoreboard_connection_TB4(1,903,3);
    `monitor_scoreboard_connection_TB4(1,904,4);
    `monitor_scoreboard_connection_TB4(1,905,5);
    `monitor_scoreboard_connection_TB4(1,906,6);
    `monitor_scoreboard_connection_TB4(1,907,7);
    `monitor_scoreboard_connection_TB4(1,908,8);
    `monitor_scoreboard_connection_TB4(1,909,9);
    `monitor_scoreboard_connection_TB4(1,910,10);
    `monitor_scoreboard_connection_TB4(1,911,11);
    `monitor_scoreboard_connection_TB4(1,912,12);
    `monitor_scoreboard_connection_TB4(1,913,13);
    `monitor_scoreboard_connection_TB4(1,914,14);
    `monitor_scoreboard_connection_TB4(1,915,15);
    `monitor_scoreboard_connection_TB4(1,916,16);
    `monitor_scoreboard_connection_TB4(1,917,17);
    `monitor_scoreboard_connection_TB4(1,918,18);
    `monitor_scoreboard_connection_TB4(1,919,19);
    `monitor_scoreboard_connection_TB4(1,920,20);
    `monitor_scoreboard_connection_TB4(1,921,21);
    `monitor_scoreboard_connection_TB4(1,922,22);
    `monitor_scoreboard_connection_TB4(1,923,23);
    `monitor_scoreboard_connection_TB4(1,924,24);
    `monitor_scoreboard_connection_TB4(1,925,25);
    `monitor_scoreboard_connection_TB4(1,926,26);
    `monitor_scoreboard_connection_TB4(1,927,27);
    `monitor_scoreboard_connection_TB4(1,928,28);
    `monitor_scoreboard_connection_TB4(1,929,29);
    `monitor_scoreboard_connection_TB4(1,930,30);
    `monitor_scoreboard_connection_TB4(1,931,31);
    `monitor_scoreboard_connection_TB4(1,932,32);
    `monitor_scoreboard_connection_TB4(1,933,33);
    `monitor_scoreboard_connection_TB4(1,934,34);
    `monitor_scoreboard_connection_TB4(1,935,35);
    `monitor_scoreboard_connection_TB4(1,936,36);
    `monitor_scoreboard_connection_TB4(1,937,37);
    `monitor_scoreboard_connection_TB4(1,938,38);
    `monitor_scoreboard_connection_TB4(1,939,39);
    `monitor_scoreboard_connection_TB4(1,940,40);
    `monitor_scoreboard_connection_TB4(1,941,41);
    `monitor_scoreboard_connection_TB4(1,942,42);
    `monitor_scoreboard_connection_TB4(1,943,43);
    `monitor_scoreboard_connection_TB4(1,944,44);
    `monitor_scoreboard_connection_TB4(1,945,45);
    `monitor_scoreboard_connection_TB4(1,946,46);
    `monitor_scoreboard_connection_TB4(1,947,47);
    `monitor_scoreboard_connection_TB4(1,948,48);
    `monitor_scoreboard_connection_TB4(1,949,49);
    `monitor_scoreboard_connection_TB4(1,950,50);
    `monitor_scoreboard_connection_TB4(1,951,51);
    `monitor_scoreboard_connection_TB4(1,952,52);
    `monitor_scoreboard_connection_TB4(1,953,53);
    `monitor_scoreboard_connection_TB4(1,954,54);
    `monitor_scoreboard_connection_TB4(1,955,55);
    `monitor_scoreboard_connection_TB4(1,956,56);
    `monitor_scoreboard_connection_TB4(1,957,57);
    `monitor_scoreboard_connection_TB4(1,958,58);
    `monitor_scoreboard_connection_TB4(1,959,59);
    `monitor_scoreboard_connection_TB4(1,960,60);
    `monitor_scoreboard_connection_TB4(1,961,61);
    `monitor_scoreboard_connection_TB4(1,962,62);
    `monitor_scoreboard_connection_TB4(1,963,63);
    `monitor_scoreboard_connection_TB4(1,964,64);
    `monitor_scoreboard_connection_TB4(1,965,65);
    `monitor_scoreboard_connection_TB4(1,966,66);
    `monitor_scoreboard_connection_TB4(1,967,67);
    `monitor_scoreboard_connection_TB4(1,968,68);
    `monitor_scoreboard_connection_TB4(1,969,69);
    `monitor_scoreboard_connection_TB4(1,970,70);
    `monitor_scoreboard_connection_TB4(1,971,71);
    `monitor_scoreboard_connection_TB4(1,972,72);
    `monitor_scoreboard_connection_TB4(1,973,73);
    `monitor_scoreboard_connection_TB4(1,974,74);
    `monitor_scoreboard_connection_TB4(1,975,75);
    `monitor_scoreboard_connection_TB4(1,976,76);
    `monitor_scoreboard_connection_TB4(1,977,77);
    `monitor_scoreboard_connection_TB4(1,978,78);
    `monitor_scoreboard_connection_TB4(1,979,79);
    `monitor_scoreboard_connection_TB4(1,980,80);
    `monitor_scoreboard_connection_TB4(1,981,81);
    `monitor_scoreboard_connection_TB4(1,982,82);
    `monitor_scoreboard_connection_TB4(1,983,83);
    `monitor_scoreboard_connection_TB4(1,984,84);
    `monitor_scoreboard_connection_TB4(1,985,85);
    `monitor_scoreboard_connection_TB4(1,986,86);
    `monitor_scoreboard_connection_TB4(1,987,87);
    `monitor_scoreboard_connection_TB4(1,988,88);
    `monitor_scoreboard_connection_TB4(1,989,89);
    `monitor_scoreboard_connection_TB4(1,990,90);
    `monitor_scoreboard_connection_TB4(1,991,91);
    `monitor_scoreboard_connection_TB4(1,992,92);
    `monitor_scoreboard_connection_TB4(1,993,93);
    `monitor_scoreboard_connection_TB4(1,994,94);
    `monitor_scoreboard_connection_TB4(1,995,95);
    `monitor_scoreboard_connection_TB4(1,996,96);
    `monitor_scoreboard_connection_TB4(1,997,97);
    `monitor_scoreboard_connection_TB4(1,998,98);
    `monitor_scoreboard_connection_TB4(1,999,99);
    `monitor_scoreboard_connection_TB4(1,1000,100);
    `monitor_scoreboard_connection_TB4(1,1001,101);
    `monitor_scoreboard_connection_TB4(1,1002,102);
    `monitor_scoreboard_connection_TB4(1,1003,103);
    `monitor_scoreboard_connection_TB4(1,1004,104);
    `monitor_scoreboard_connection_TB4(1,1005,105);
    `monitor_scoreboard_connection_TB4(1,1006,106);
    `monitor_scoreboard_connection_TB4(1,1007,107);
    `monitor_scoreboard_connection_TB4(1,1008,108);
    `monitor_scoreboard_connection_TB4(1,1009,109);
    `monitor_scoreboard_connection_TB4(1,1010,110);
    `monitor_scoreboard_connection_TB4(1,1011,111);
    `monitor_scoreboard_connection_TB4(1,1012,112);
    `monitor_scoreboard_connection_TB4(1,1013,113);
    `monitor_scoreboard_connection_TB4(1,1014,114);
    `monitor_scoreboard_connection_TB4(1,1015,115);
    `monitor_scoreboard_connection_TB4(1,1016,116);
    `monitor_scoreboard_connection_TB4(1,1017,117);
    `monitor_scoreboard_connection_TB4(1,1018,118);
    `monitor_scoreboard_connection_TB4(1,1019,119);
    `monitor_scoreboard_connection_TB4(1,1020,120);
    `monitor_scoreboard_connection_TB4(1,1021,121);
    `monitor_scoreboard_connection_TB4(1,1022,122);
    `monitor_scoreboard_connection_TB4(1,1023,123);
    `monitor_scoreboard_connection_TB4(1,1024,124);
    `monitor_scoreboard_connection_TB4(1,1025,125);
    `monitor_scoreboard_connection_TB4(1,1026,126);
    `monitor_scoreboard_connection_TB4(1,1027,127);
    `monitor_scoreboard_connection_TB4(1,1028,128);
    `monitor_scoreboard_connection_TB4(1,1029,129);
    `monitor_scoreboard_connection_TB4(1,1030,130);
    `monitor_scoreboard_connection_TB4(1,1031,131);
    `monitor_scoreboard_connection_TB4(1,1032,132);
    `monitor_scoreboard_connection_TB4(1,1033,133);
    `monitor_scoreboard_connection_TB4(1,1034,134);
    `monitor_scoreboard_connection_TB4(1,1035,135);
    `monitor_scoreboard_connection_TB4(1,1036,136);
    `monitor_scoreboard_connection_TB4(1,1037,137);
    `monitor_scoreboard_connection_TB4(1,1038,138);
    `monitor_scoreboard_connection_TB4(1,1039,139);
    `monitor_scoreboard_connection_TB4(1,1040,140);
    `monitor_scoreboard_connection_TB4(1,1041,141);
    `monitor_scoreboard_connection_TB4(1,1042,142);
    `monitor_scoreboard_connection_TB4(1,1043,143);
    `monitor_scoreboard_connection_TB4(1,1044,144);
    `monitor_scoreboard_connection_TB4(1,1045,145);
    `monitor_scoreboard_connection_TB4(1,1046,146);
    `monitor_scoreboard_connection_TB4(1,1047,147);
    `monitor_scoreboard_connection_TB4(1,1048,148);
    `monitor_scoreboard_connection_TB4(1,1049,149);
    `monitor_scoreboard_connection_TB4(1,1050,150);
    `monitor_scoreboard_connection_TB4(1,1051,151);
    `monitor_scoreboard_connection_TB4(1,1052,152);
    `monitor_scoreboard_connection_TB4(1,1053,153);
    `monitor_scoreboard_connection_TB4(1,1054,154);
    `monitor_scoreboard_connection_TB4(1,1055,155);
    `monitor_scoreboard_connection_TB4(1,1056,156);
    `monitor_scoreboard_connection_TB4(1,1057,157);
    `monitor_scoreboard_connection_TB4(1,1058,158);
    `monitor_scoreboard_connection_TB4(1,1059,159);
    `monitor_scoreboard_connection_TB4(1,1060,160);
    `monitor_scoreboard_connection_TB4(1,1061,161);
    `monitor_scoreboard_connection_TB4(1,1062,162);
    `monitor_scoreboard_connection_TB4(1,1063,163);
    `monitor_scoreboard_connection_TB4(1,1064,164);
    `monitor_scoreboard_connection_TB4(1,1065,165);
    `monitor_scoreboard_connection_TB4(1,1066,166);
    `monitor_scoreboard_connection_TB4(1,1067,167);
    `monitor_scoreboard_connection_TB4(1,1068,168);
    `monitor_scoreboard_connection_TB4(1,1069,169);
    `monitor_scoreboard_connection_TB4(1,1070,170);
    `monitor_scoreboard_connection_TB4(1,1071,171);
    `monitor_scoreboard_connection_TB4(1,1072,172);
    `monitor_scoreboard_connection_TB4(1,1073,173);
    `monitor_scoreboard_connection_TB4(1,1074,174);
    `monitor_scoreboard_connection_TB4(1,1075,175);
    `monitor_scoreboard_connection_TB4(1,1076,176);
    `monitor_scoreboard_connection_TB4(1,1077,177);
    `monitor_scoreboard_connection_TB4(1,1078,178);
    `monitor_scoreboard_connection_TB4(1,1079,179);
    `monitor_scoreboard_connection_TB4(1,1080,180);
    `monitor_scoreboard_connection_TB4(1,1081,181);
    `monitor_scoreboard_connection_TB4(1,1082,182);
    `monitor_scoreboard_connection_TB4(1,1083,183);
    `monitor_scoreboard_connection_TB4(1,1084,184);
    `monitor_scoreboard_connection_TB4(1,1085,185);
    `monitor_scoreboard_connection_TB4(1,1086,186);
    `monitor_scoreboard_connection_TB4(1,1087,187);
    `monitor_scoreboard_connection_TB4(1,1088,188);
    `monitor_scoreboard_connection_TB4(1,1089,189);
    `monitor_scoreboard_connection_TB4(1,1090,190);
    `monitor_scoreboard_connection_TB4(1,1091,191);
    `monitor_scoreboard_connection_TB4(1,1092,192);
    `monitor_scoreboard_connection_TB4(1,1093,193);
    `monitor_scoreboard_connection_TB4(1,1094,194);
    `monitor_scoreboard_connection_TB4(1,1095,195);
    `monitor_scoreboard_connection_TB4(1,1096,196);
    `monitor_scoreboard_connection_TB4(1,1097,197);
    `monitor_scoreboard_connection_TB4(1,1098,198);
    `monitor_scoreboard_connection_TB4(1,1099,199);
    `monitor_scoreboard_connection_TB4(1,1100,200);
    `monitor_scoreboard_connection_TB4(1,1101,201);
    `monitor_scoreboard_connection_TB4(1,1102,202);
    `monitor_scoreboard_connection_TB4(1,1103,203);
    `monitor_scoreboard_connection_TB4(1,1104,204);
    `monitor_scoreboard_connection_TB4(1,1105,205);
    `monitor_scoreboard_connection_TB4(1,1106,206);
    `monitor_scoreboard_connection_TB4(1,1107,207);
    `monitor_scoreboard_connection_TB4(1,1108,208);
    `monitor_scoreboard_connection_TB4(1,1109,209);
    `monitor_scoreboard_connection_TB4(1,1110,210);
    `monitor_scoreboard_connection_TB4(1,1111,211);
    `monitor_scoreboard_connection_TB4(1,1112,212);
    `monitor_scoreboard_connection_TB4(1,1113,213);
    `monitor_scoreboard_connection_TB4(1,1114,214);
    `monitor_scoreboard_connection_TB4(1,1115,215);
    `monitor_scoreboard_connection_TB4(1,1116,216);
    `monitor_scoreboard_connection_TB4(1,1117,217);
    `monitor_scoreboard_connection_TB4(1,1118,218);
    `monitor_scoreboard_connection_TB4(1,1119,219);
    `monitor_scoreboard_connection_TB4(1,1120,220);
    `monitor_scoreboard_connection_TB4(1,1121,221);
    `monitor_scoreboard_connection_TB4(1,1122,222);
    `monitor_scoreboard_connection_TB4(1,1123,223);
    `monitor_scoreboard_connection_TB4(1,1124,224);
    `monitor_scoreboard_connection_TB4(1,1125,225);
    `monitor_scoreboard_connection_TB4(1,1126,226);
    `monitor_scoreboard_connection_TB4(1,1127,227);
    `monitor_scoreboard_connection_TB4(1,1128,228);
    `monitor_scoreboard_connection_TB4(1,1129,229);
    `monitor_scoreboard_connection_TB4(1,1130,230);
    `monitor_scoreboard_connection_TB4(1,1131,231);
    `monitor_scoreboard_connection_TB4(1,1132,232);
    `monitor_scoreboard_connection_TB4(1,1133,233);
    `monitor_scoreboard_connection_TB4(1,1134,234);
    `monitor_scoreboard_connection_TB4(1,1135,235);
    `monitor_scoreboard_connection_TB4(1,1136,236);
    `monitor_scoreboard_connection_TB4(1,1137,237);
    `monitor_scoreboard_connection_TB4(1,1138,238);
    `monitor_scoreboard_connection_TB4(1,1139,239);
    `monitor_scoreboard_connection_TB4(1,1140,240);
    `monitor_scoreboard_connection_TB4(1,1141,241);
    `monitor_scoreboard_connection_TB4(1,1142,242);
    `monitor_scoreboard_connection_TB4(1,1143,243);
    `monitor_scoreboard_connection_TB4(1,1144,244);
    `monitor_scoreboard_connection_TB4(1,1145,245);
    `monitor_scoreboard_connection_TB4(1,1146,246);
    `monitor_scoreboard_connection_TB4(1,1147,247);
    `monitor_scoreboard_connection_TB4(1,1148,248);
    `monitor_scoreboard_connection_TB4(1,1149,249);
    `monitor_scoreboard_connection_TB4(1,1150,250);
    `monitor_scoreboard_connection_TB4(1,1151,251);
    `monitor_scoreboard_connection_TB4(1,1152,252);
    `monitor_scoreboard_connection_TB4(1,1153,253);
    `monitor_scoreboard_connection_TB4(1,1154,254);
    `monitor_scoreboard_connection_TB4(1,1155,255);
    `monitor_scoreboard_connection_TB4(1,1156,256);
    `monitor_scoreboard_connection_TB4(1,1157,257);
    `monitor_scoreboard_connection_TB4(1,1158,258);
    `monitor_scoreboard_connection_TB4(1,1159,259);
    `monitor_scoreboard_connection_TB4(1,1160,260);
    `monitor_scoreboard_connection_TB4(1,1161,261);
    `monitor_scoreboard_connection_TB4(1,1162,262);
    `monitor_scoreboard_connection_TB4(1,1163,263);
    `monitor_scoreboard_connection_TB4(1,1164,264);
    `monitor_scoreboard_connection_TB4(1,1165,265);
    `monitor_scoreboard_connection_TB4(1,1166,266);
    `monitor_scoreboard_connection_TB4(1,1167,267);
    `monitor_scoreboard_connection_TB4(1,1168,268);
    `monitor_scoreboard_connection_TB4(1,1169,269);
    `monitor_scoreboard_connection_TB4(1,1170,270);
    `monitor_scoreboard_connection_TB4(1,1171,271);
    `monitor_scoreboard_connection_TB4(1,1172,272);
    `monitor_scoreboard_connection_TB4(1,1173,273);
    `monitor_scoreboard_connection_TB4(1,1174,274);
    `monitor_scoreboard_connection_TB4(1,1175,275);
    `monitor_scoreboard_connection_TB4(1,1176,276);
    `monitor_scoreboard_connection_TB4(1,1177,277);
    `monitor_scoreboard_connection_TB4(1,1178,278);
    `monitor_scoreboard_connection_TB4(1,1179,279);
    `monitor_scoreboard_connection_TB4(1,1180,280);
    `monitor_scoreboard_connection_TB4(1,1181,281);
    `monitor_scoreboard_connection_TB4(1,1182,282);
    `monitor_scoreboard_connection_TB4(1,1183,283);
    `monitor_scoreboard_connection_TB4(1,1184,284);
    `monitor_scoreboard_connection_TB4(1,1185,285);
    `monitor_scoreboard_connection_TB4(1,1186,286);
    `monitor_scoreboard_connection_TB4(1,1187,287);
    `monitor_scoreboard_connection_TB4(1,1188,288);
    `monitor_scoreboard_connection_TB4(1,1189,289);
    `monitor_scoreboard_connection_TB4(1,1190,290);
    `monitor_scoreboard_connection_TB4(1,1191,291);
    `monitor_scoreboard_connection_TB4(1,1192,292);
    `monitor_scoreboard_connection_TB4(1,1193,293);
    `monitor_scoreboard_connection_TB4(1,1194,294);
    `monitor_scoreboard_connection_TB4(1,1195,295);
    `monitor_scoreboard_connection_TB4(1,1196,296);
    `monitor_scoreboard_connection_TB4(1,1197,297);
    `monitor_scoreboard_connection_TB4(1,1198,298);
    `monitor_scoreboard_connection_TB4(1,1199,299);
    `monitor_scoreboard_connection_TB4(1,1200,300);
    `monitor_scoreboard_connection_TB4(1,1201,301);
    `monitor_scoreboard_connection_TB4(1,1202,302);
    `monitor_scoreboard_connection_TB4(1,1203,303);
    `monitor_scoreboard_connection_TB4(1,1204,304);
    `monitor_scoreboard_connection_TB4(1,1205,305);
    `monitor_scoreboard_connection_TB4(1,1206,306);
    `monitor_scoreboard_connection_TB4(1,1207,307);
    `monitor_scoreboard_connection_TB4(1,1208,308);
    `monitor_scoreboard_connection_TB4(1,1209,309);
    `monitor_scoreboard_connection_TB4(1,1210,310);
    `monitor_scoreboard_connection_TB4(1,1211,311);
    `monitor_scoreboard_connection_TB4(1,1212,312);
    `monitor_scoreboard_connection_TB4(1,1213,313);
    `monitor_scoreboard_connection_TB4(1,1214,314);
    `monitor_scoreboard_connection_TB4(1,1215,315);
    `monitor_scoreboard_connection_TB4(1,1216,316);
    `monitor_scoreboard_connection_TB4(1,1217,317);
    `monitor_scoreboard_connection_TB4(1,1218,318);
    `monitor_scoreboard_connection_TB4(1,1219,319);
    `monitor_scoreboard_connection_TB4(1,1220,320);
    `monitor_scoreboard_connection_TB4(1,1221,321);
    `monitor_scoreboard_connection_TB4(1,1222,322);
    `monitor_scoreboard_connection_TB4(1,1223,323);
    `monitor_scoreboard_connection_TB4(1,1224,324);
    `monitor_scoreboard_connection_TB4(1,1225,325);
    `monitor_scoreboard_connection_TB4(1,1226,326);
    `monitor_scoreboard_connection_TB4(1,1227,327);
    `monitor_scoreboard_connection_TB4(1,1228,328);
    `monitor_scoreboard_connection_TB4(1,1229,329);
    `monitor_scoreboard_connection_TB4(1,1230,330);
    `monitor_scoreboard_connection_TB4(1,1231,331);
    `monitor_scoreboard_connection_TB4(1,1232,332);
    `monitor_scoreboard_connection_TB4(1,1233,333);
    `monitor_scoreboard_connection_TB4(1,1234,334);
    `monitor_scoreboard_connection_TB4(1,1235,335);
    `monitor_scoreboard_connection_TB4(1,1236,336);
    `monitor_scoreboard_connection_TB4(1,1237,337);
    `monitor_scoreboard_connection_TB4(1,1238,338);
    `monitor_scoreboard_connection_TB4(1,1239,339);
    `monitor_scoreboard_connection_TB4(1,1240,340);
    `monitor_scoreboard_connection_TB4(1,1241,341);
    `monitor_scoreboard_connection_TB4(1,1242,342);
    `monitor_scoreboard_connection_TB4(1,1243,343);
    `monitor_scoreboard_connection_TB4(1,1244,344);
    `monitor_scoreboard_connection_TB4(1,1245,345);
    `monitor_scoreboard_connection_TB4(1,1246,346);
    `monitor_scoreboard_connection_TB4(1,1247,347);
    `monitor_scoreboard_connection_TB4(1,1248,348);
    `monitor_scoreboard_connection_TB4(1,1249,349);
    `monitor_scoreboard_connection_TB4(1,1250,350);
    `monitor_scoreboard_connection_TB4(1,1251,351);
    `monitor_scoreboard_connection_TB4(1,1252,352);
    `monitor_scoreboard_connection_TB4(1,1253,353);
    `monitor_scoreboard_connection_TB4(1,1254,354);
    `monitor_scoreboard_connection_TB4(1,1255,355);
    `monitor_scoreboard_connection_TB4(1,1256,356);
    `monitor_scoreboard_connection_TB4(1,1257,357);
    `monitor_scoreboard_connection_TB4(1,1258,358);
    `monitor_scoreboard_connection_TB4(1,1259,359);
    `monitor_scoreboard_connection_TB4(1,1260,360);
    `monitor_scoreboard_connection_TB4(1,1261,361);
    `monitor_scoreboard_connection_TB4(1,1262,362);
    `monitor_scoreboard_connection_TB4(1,1263,363);
    `monitor_scoreboard_connection_TB4(1,1264,364);
    `monitor_scoreboard_connection_TB4(1,1265,365);
    `monitor_scoreboard_connection_TB4(1,1266,366);
    `monitor_scoreboard_connection_TB4(1,1267,367);
    `monitor_scoreboard_connection_TB4(1,1268,368);
    `monitor_scoreboard_connection_TB4(1,1269,369);
    `monitor_scoreboard_connection_TB4(1,1270,370);
    `monitor_scoreboard_connection_TB4(1,1271,371);
    `monitor_scoreboard_connection_TB4(1,1272,372);
    `monitor_scoreboard_connection_TB4(1,1273,373);
    `monitor_scoreboard_connection_TB4(1,1274,374);
    `monitor_scoreboard_connection_TB4(1,1275,375);
    `monitor_scoreboard_connection_TB4(1,1276,376);
    `monitor_scoreboard_connection_TB4(1,1277,377);
    `monitor_scoreboard_connection_TB4(1,1278,378);
    `monitor_scoreboard_connection_TB4(1,1279,379);
    `monitor_scoreboard_connection_TB4(1,1280,380);
    `monitor_scoreboard_connection_TB4(1,1281,381);
    `monitor_scoreboard_connection_TB4(1,1282,382);
    `monitor_scoreboard_connection_TB4(1,1283,383);
    `monitor_scoreboard_connection_TB4(1,1284,384);
    `monitor_scoreboard_connection_TB4(1,1285,385);
    `monitor_scoreboard_connection_TB4(1,1286,386);
    `monitor_scoreboard_connection_TB4(1,1287,387);
    `monitor_scoreboard_connection_TB4(1,1288,388);
    `monitor_scoreboard_connection_TB4(1,1289,389);
    `monitor_scoreboard_connection_TB4(1,1290,390);
    `monitor_scoreboard_connection_TB4(1,1291,391);
    `monitor_scoreboard_connection_TB4(1,1292,392);
    `monitor_scoreboard_connection_TB4(1,1293,393);
    `monitor_scoreboard_connection_TB4(1,1294,394);
    `monitor_scoreboard_connection_TB4(1,1295,395);
    `monitor_scoreboard_connection_TB4(1,1296,396);
    `monitor_scoreboard_connection_TB4(1,1297,397);
    `monitor_scoreboard_connection_TB4(1,1298,398);
    `monitor_scoreboard_connection_TB4(1,1299,399);
    `monitor_scoreboard_connection_TB4(1,1300,400);
    `monitor_scoreboard_connection_TB4(1,1301,401);
    `monitor_scoreboard_connection_TB4(1,1302,402);
    `monitor_scoreboard_connection_TB4(1,1303,403);
    `monitor_scoreboard_connection_TB4(1,1304,404);
    `monitor_scoreboard_connection_TB4(1,1305,405);
    `monitor_scoreboard_connection_TB4(1,1306,406);
    `monitor_scoreboard_connection_TB4(1,1307,407);
    `monitor_scoreboard_connection_TB4(1,1308,408);
    `monitor_scoreboard_connection_TB4(1,1309,409);
    `monitor_scoreboard_connection_TB4(1,1310,410);
    `monitor_scoreboard_connection_TB4(1,1311,411);
    `monitor_scoreboard_connection_TB4(1,1312,412);
    `monitor_scoreboard_connection_TB4(1,1313,413);
    `monitor_scoreboard_connection_TB4(1,1314,414);
    `monitor_scoreboard_connection_TB4(1,1315,415);
    `monitor_scoreboard_connection_TB4(1,1316,416);
    `monitor_scoreboard_connection_TB4(1,1317,417);
    `monitor_scoreboard_connection_TB4(1,1318,418);
    `monitor_scoreboard_connection_TB4(1,1319,419);
    `monitor_scoreboard_connection_TB4(1,1320,420);
    `monitor_scoreboard_connection_TB4(1,1321,421);
    `monitor_scoreboard_connection_TB4(1,1322,422);
    `monitor_scoreboard_connection_TB4(1,1323,423);
    `monitor_scoreboard_connection_TB4(1,1324,424);
    `monitor_scoreboard_connection_TB4(1,1325,425);
    `monitor_scoreboard_connection_TB4(1,1326,426);
    `monitor_scoreboard_connection_TB4(1,1327,427);
    `monitor_scoreboard_connection_TB4(1,1328,428);
    `monitor_scoreboard_connection_TB4(1,1329,429);
    `monitor_scoreboard_connection_TB4(1,1330,430);
    `monitor_scoreboard_connection_TB4(1,1331,431);
    `monitor_scoreboard_connection_TB4(1,1332,432);
    `monitor_scoreboard_connection_TB4(1,1333,433);
    `monitor_scoreboard_connection_TB4(1,1334,434);
    `monitor_scoreboard_connection_TB4(1,1335,435);
    `monitor_scoreboard_connection_TB4(1,1336,436);
    `monitor_scoreboard_connection_TB4(1,1337,437);
    `monitor_scoreboard_connection_TB4(1,1338,438);
    `monitor_scoreboard_connection_TB4(1,1339,439);
    `monitor_scoreboard_connection_TB4(1,1340,440);
    `monitor_scoreboard_connection_TB4(1,1341,441);
    `monitor_scoreboard_connection_TB4(1,1342,442);
    `monitor_scoreboard_connection_TB4(1,1343,443);
    `monitor_scoreboard_connection_TB4(1,1344,444);
    `monitor_scoreboard_connection_TB4(1,1345,445);
    `monitor_scoreboard_connection_TB4(1,1346,446);
    `monitor_scoreboard_connection_TB4(1,1347,447);
    `monitor_scoreboard_connection_TB4(1,1348,448);
    `monitor_scoreboard_connection_TB4(1,1349,449);
    `monitor_scoreboard_connection_TB4(2,1350,0);
    `monitor_scoreboard_connection_TB4(2,1351,1);
    `monitor_scoreboard_connection_TB4(2,1352,2);
    `monitor_scoreboard_connection_TB4(2,1353,3);
    `monitor_scoreboard_connection_TB4(2,1354,4);
    `monitor_scoreboard_connection_TB4(2,1355,5);
    `monitor_scoreboard_connection_TB4(2,1356,6);
    `monitor_scoreboard_connection_TB4(2,1357,7);
    `monitor_scoreboard_connection_TB4(2,1358,8);
    `monitor_scoreboard_connection_TB4(2,1359,9);
    `monitor_scoreboard_connection_TB4(2,1360,10);
    `monitor_scoreboard_connection_TB4(2,1361,11);
    `monitor_scoreboard_connection_TB4(2,1362,12);
    `monitor_scoreboard_connection_TB4(2,1363,13);
    `monitor_scoreboard_connection_TB4(2,1364,14);
    `monitor_scoreboard_connection_TB4(2,1365,15);
    `monitor_scoreboard_connection_TB4(2,1366,16);
    `monitor_scoreboard_connection_TB4(2,1367,17);
    `monitor_scoreboard_connection_TB4(2,1368,18);
    `monitor_scoreboard_connection_TB4(2,1369,19);
    `monitor_scoreboard_connection_TB4(2,1370,20);
    `monitor_scoreboard_connection_TB4(2,1371,21);
    `monitor_scoreboard_connection_TB4(2,1372,22);
    `monitor_scoreboard_connection_TB4(2,1373,23);
    `monitor_scoreboard_connection_TB4(2,1374,24);
    `monitor_scoreboard_connection_TB4(2,1375,25);
    `monitor_scoreboard_connection_TB4(2,1376,26);
    `monitor_scoreboard_connection_TB4(2,1377,27);
    `monitor_scoreboard_connection_TB4(2,1378,28);
    `monitor_scoreboard_connection_TB4(2,1379,29);
    `monitor_scoreboard_connection_TB4(2,1380,30);
    `monitor_scoreboard_connection_TB4(2,1381,31);
    `monitor_scoreboard_connection_TB4(2,1382,32);
    `monitor_scoreboard_connection_TB4(2,1383,33);
    `monitor_scoreboard_connection_TB4(2,1384,34);
    `monitor_scoreboard_connection_TB4(2,1385,35);
    `monitor_scoreboard_connection_TB4(2,1386,36);
    `monitor_scoreboard_connection_TB4(2,1387,37);
    `monitor_scoreboard_connection_TB4(2,1388,38);
    `monitor_scoreboard_connection_TB4(2,1389,39);
    `monitor_scoreboard_connection_TB4(2,1390,40);
    `monitor_scoreboard_connection_TB4(2,1391,41);
    `monitor_scoreboard_connection_TB4(2,1392,42);
    `monitor_scoreboard_connection_TB4(2,1393,43);
    `monitor_scoreboard_connection_TB4(2,1394,44);
    `monitor_scoreboard_connection_TB4(2,1395,45);
    `monitor_scoreboard_connection_TB4(2,1396,46);
    `monitor_scoreboard_connection_TB4(2,1397,47);
    `monitor_scoreboard_connection_TB4(2,1398,48);
    `monitor_scoreboard_connection_TB4(2,1399,49);
    `monitor_scoreboard_connection_TB4(2,1400,50);
    `monitor_scoreboard_connection_TB4(2,1401,51);
    `monitor_scoreboard_connection_TB4(2,1402,52);
    `monitor_scoreboard_connection_TB4(2,1403,53);
    `monitor_scoreboard_connection_TB4(2,1404,54);
    `monitor_scoreboard_connection_TB4(2,1405,55);
    `monitor_scoreboard_connection_TB4(2,1406,56);
    `monitor_scoreboard_connection_TB4(2,1407,57);
    `monitor_scoreboard_connection_TB4(2,1408,58);
    `monitor_scoreboard_connection_TB4(2,1409,59);
    `monitor_scoreboard_connection_TB4(2,1410,60);
    `monitor_scoreboard_connection_TB4(2,1411,61);
    `monitor_scoreboard_connection_TB4(2,1412,62);
    `monitor_scoreboard_connection_TB4(2,1413,63);
    `monitor_scoreboard_connection_TB4(2,1414,64);
    `monitor_scoreboard_connection_TB4(2,1415,65);
    `monitor_scoreboard_connection_TB4(2,1416,66);
    `monitor_scoreboard_connection_TB4(2,1417,67);
    `monitor_scoreboard_connection_TB4(2,1418,68);
    `monitor_scoreboard_connection_TB4(2,1419,69);
    `monitor_scoreboard_connection_TB4(2,1420,70);
    `monitor_scoreboard_connection_TB4(2,1421,71);
    `monitor_scoreboard_connection_TB4(2,1422,72);
    `monitor_scoreboard_connection_TB4(2,1423,73);
    `monitor_scoreboard_connection_TB4(2,1424,74);
    `monitor_scoreboard_connection_TB4(2,1425,75);
    `monitor_scoreboard_connection_TB4(2,1426,76);
    `monitor_scoreboard_connection_TB4(2,1427,77);
    `monitor_scoreboard_connection_TB4(2,1428,78);
    `monitor_scoreboard_connection_TB4(2,1429,79);
    `monitor_scoreboard_connection_TB4(2,1430,80);
    `monitor_scoreboard_connection_TB4(2,1431,81);
    `monitor_scoreboard_connection_TB4(2,1432,82);
    `monitor_scoreboard_connection_TB4(2,1433,83);
    `monitor_scoreboard_connection_TB4(2,1434,84);
    `monitor_scoreboard_connection_TB4(2,1435,85);
    `monitor_scoreboard_connection_TB4(2,1436,86);
    `monitor_scoreboard_connection_TB4(2,1437,87);
    `monitor_scoreboard_connection_TB4(2,1438,88);
    `monitor_scoreboard_connection_TB4(2,1439,89);
    `monitor_scoreboard_connection_TB4(2,1440,90);
    `monitor_scoreboard_connection_TB4(2,1441,91);
    `monitor_scoreboard_connection_TB4(2,1442,92);
    `monitor_scoreboard_connection_TB4(2,1443,93);
    `monitor_scoreboard_connection_TB4(2,1444,94);
    `monitor_scoreboard_connection_TB4(2,1445,95);
    `monitor_scoreboard_connection_TB4(2,1446,96);
    `monitor_scoreboard_connection_TB4(2,1447,97);
    `monitor_scoreboard_connection_TB4(2,1448,98);
    `monitor_scoreboard_connection_TB4(2,1449,99);
    `monitor_scoreboard_connection_TB4(2,1450,100);
    `monitor_scoreboard_connection_TB4(2,1451,101);
    `monitor_scoreboard_connection_TB4(2,1452,102);
    `monitor_scoreboard_connection_TB4(2,1453,103);
    `monitor_scoreboard_connection_TB4(2,1454,104);
    `monitor_scoreboard_connection_TB4(2,1455,105);
    `monitor_scoreboard_connection_TB4(2,1456,106);
    `monitor_scoreboard_connection_TB4(2,1457,107);
    `monitor_scoreboard_connection_TB4(2,1458,108);
    `monitor_scoreboard_connection_TB4(2,1459,109);
    `monitor_scoreboard_connection_TB4(2,1460,110);
    `monitor_scoreboard_connection_TB4(2,1461,111);
    `monitor_scoreboard_connection_TB4(2,1462,112);
    `monitor_scoreboard_connection_TB4(2,1463,113);
    `monitor_scoreboard_connection_TB4(2,1464,114);
    `monitor_scoreboard_connection_TB4(2,1465,115);
    `monitor_scoreboard_connection_TB4(2,1466,116);
    `monitor_scoreboard_connection_TB4(2,1467,117);
    `monitor_scoreboard_connection_TB4(2,1468,118);
    `monitor_scoreboard_connection_TB4(2,1469,119);
    `monitor_scoreboard_connection_TB4(2,1470,120);
    `monitor_scoreboard_connection_TB4(2,1471,121);
    `monitor_scoreboard_connection_TB4(2,1472,122);
    `monitor_scoreboard_connection_TB4(2,1473,123);
    `monitor_scoreboard_connection_TB4(2,1474,124);
    `monitor_scoreboard_connection_TB4(2,1475,125);
    `monitor_scoreboard_connection_TB4(2,1476,126);
    `monitor_scoreboard_connection_TB4(2,1477,127);
    `monitor_scoreboard_connection_TB4(2,1478,128);
    `monitor_scoreboard_connection_TB4(2,1479,129);
    `monitor_scoreboard_connection_TB4(2,1480,130);
    `monitor_scoreboard_connection_TB4(2,1481,131);
    `monitor_scoreboard_connection_TB4(2,1482,132);
    `monitor_scoreboard_connection_TB4(2,1483,133);
    `monitor_scoreboard_connection_TB4(2,1484,134);
    `monitor_scoreboard_connection_TB4(2,1485,135);
    `monitor_scoreboard_connection_TB4(2,1486,136);
    `monitor_scoreboard_connection_TB4(2,1487,137);
    `monitor_scoreboard_connection_TB4(2,1488,138);
    `monitor_scoreboard_connection_TB4(2,1489,139);
    `monitor_scoreboard_connection_TB4(2,1490,140);
    `monitor_scoreboard_connection_TB4(2,1491,141);
    `monitor_scoreboard_connection_TB4(2,1492,142);
    `monitor_scoreboard_connection_TB4(2,1493,143);
    `monitor_scoreboard_connection_TB4(2,1494,144);
    `monitor_scoreboard_connection_TB4(2,1495,145);
    `monitor_scoreboard_connection_TB4(2,1496,146);
    `monitor_scoreboard_connection_TB4(2,1497,147);
    `monitor_scoreboard_connection_TB4(2,1498,148);
    `monitor_scoreboard_connection_TB4(2,1499,149);
    `monitor_scoreboard_connection_TB4(2,1500,150);
    `monitor_scoreboard_connection_TB4(2,1501,151);
    `monitor_scoreboard_connection_TB4(2,1502,152);
    `monitor_scoreboard_connection_TB4(2,1503,153);
    `monitor_scoreboard_connection_TB4(2,1504,154);
    `monitor_scoreboard_connection_TB4(2,1505,155);
    `monitor_scoreboard_connection_TB4(2,1506,156);
    `monitor_scoreboard_connection_TB4(2,1507,157);
    `monitor_scoreboard_connection_TB4(2,1508,158);
    `monitor_scoreboard_connection_TB4(2,1509,159);
    `monitor_scoreboard_connection_TB4(2,1510,160);
    `monitor_scoreboard_connection_TB4(2,1511,161);
    `monitor_scoreboard_connection_TB4(2,1512,162);
    `monitor_scoreboard_connection_TB4(2,1513,163);
    `monitor_scoreboard_connection_TB4(2,1514,164);
    `monitor_scoreboard_connection_TB4(2,1515,165);
    `monitor_scoreboard_connection_TB4(2,1516,166);
    `monitor_scoreboard_connection_TB4(2,1517,167);
    `monitor_scoreboard_connection_TB4(2,1518,168);
    `monitor_scoreboard_connection_TB4(2,1519,169);
    `monitor_scoreboard_connection_TB4(2,1520,170);
    `monitor_scoreboard_connection_TB4(2,1521,171);
    `monitor_scoreboard_connection_TB4(2,1522,172);
    `monitor_scoreboard_connection_TB4(2,1523,173);
    `monitor_scoreboard_connection_TB4(2,1524,174);
    `monitor_scoreboard_connection_TB4(2,1525,175);
    `monitor_scoreboard_connection_TB4(2,1526,176);
    `monitor_scoreboard_connection_TB4(2,1527,177);
    `monitor_scoreboard_connection_TB4(2,1528,178);
    `monitor_scoreboard_connection_TB4(2,1529,179);
    `monitor_scoreboard_connection_TB4(2,1530,180);
    `monitor_scoreboard_connection_TB4(2,1531,181);
    `monitor_scoreboard_connection_TB4(2,1532,182);
    `monitor_scoreboard_connection_TB4(2,1533,183);
    `monitor_scoreboard_connection_TB4(2,1534,184);
    `monitor_scoreboard_connection_TB4(2,1535,185);
    `monitor_scoreboard_connection_TB4(2,1536,186);
    `monitor_scoreboard_connection_TB4(2,1537,187);
    `monitor_scoreboard_connection_TB4(2,1538,188);
    `monitor_scoreboard_connection_TB4(2,1539,189);
    `monitor_scoreboard_connection_TB4(2,1540,190);
    `monitor_scoreboard_connection_TB4(2,1541,191);
    `monitor_scoreboard_connection_TB4(2,1542,192);
    `monitor_scoreboard_connection_TB4(2,1543,193);
    `monitor_scoreboard_connection_TB4(2,1544,194);
    `monitor_scoreboard_connection_TB4(2,1545,195);
    `monitor_scoreboard_connection_TB4(2,1546,196);
    `monitor_scoreboard_connection_TB4(2,1547,197);
    `monitor_scoreboard_connection_TB4(2,1548,198);
    `monitor_scoreboard_connection_TB4(2,1549,199);
    `monitor_scoreboard_connection_TB4(2,1550,200);
    `monitor_scoreboard_connection_TB4(2,1551,201);
    `monitor_scoreboard_connection_TB4(2,1552,202);
    `monitor_scoreboard_connection_TB4(2,1553,203);
    `monitor_scoreboard_connection_TB4(2,1554,204);
    `monitor_scoreboard_connection_TB4(2,1555,205);
    `monitor_scoreboard_connection_TB4(2,1556,206);
    `monitor_scoreboard_connection_TB4(2,1557,207);
    `monitor_scoreboard_connection_TB4(2,1558,208);
    `monitor_scoreboard_connection_TB4(2,1559,209);
    `monitor_scoreboard_connection_TB4(2,1560,210);
    `monitor_scoreboard_connection_TB4(2,1561,211);
    `monitor_scoreboard_connection_TB4(2,1562,212);
    `monitor_scoreboard_connection_TB4(2,1563,213);
    `monitor_scoreboard_connection_TB4(2,1564,214);
    `monitor_scoreboard_connection_TB4(2,1565,215);
    `monitor_scoreboard_connection_TB4(2,1566,216);
    `monitor_scoreboard_connection_TB4(2,1567,217);
    `monitor_scoreboard_connection_TB4(2,1568,218);
    `monitor_scoreboard_connection_TB4(2,1569,219);
    `monitor_scoreboard_connection_TB4(2,1570,220);
    `monitor_scoreboard_connection_TB4(2,1571,221);
    `monitor_scoreboard_connection_TB4(2,1572,222);
    `monitor_scoreboard_connection_TB4(2,1573,223);
    `monitor_scoreboard_connection_TB4(2,1574,224);
    `monitor_scoreboard_connection_TB4(2,1575,225);
    `monitor_scoreboard_connection_TB4(2,1576,226);
    `monitor_scoreboard_connection_TB4(2,1577,227);
    `monitor_scoreboard_connection_TB4(2,1578,228);
    `monitor_scoreboard_connection_TB4(2,1579,229);
    `monitor_scoreboard_connection_TB4(2,1580,230);
    `monitor_scoreboard_connection_TB4(2,1581,231);
    `monitor_scoreboard_connection_TB4(2,1582,232);
    `monitor_scoreboard_connection_TB4(2,1583,233);
    `monitor_scoreboard_connection_TB4(2,1584,234);
    `monitor_scoreboard_connection_TB4(2,1585,235);
    `monitor_scoreboard_connection_TB4(2,1586,236);
    `monitor_scoreboard_connection_TB4(2,1587,237);
    `monitor_scoreboard_connection_TB4(2,1588,238);
    `monitor_scoreboard_connection_TB4(2,1589,239);
    `monitor_scoreboard_connection_TB4(2,1590,240);
    `monitor_scoreboard_connection_TB4(2,1591,241);
    `monitor_scoreboard_connection_TB4(2,1592,242);
    `monitor_scoreboard_connection_TB4(2,1593,243);
    `monitor_scoreboard_connection_TB4(2,1594,244);
    `monitor_scoreboard_connection_TB4(2,1595,245);
    `monitor_scoreboard_connection_TB4(2,1596,246);
    `monitor_scoreboard_connection_TB4(2,1597,247);
    `monitor_scoreboard_connection_TB4(2,1598,248);
    `monitor_scoreboard_connection_TB4(2,1599,249);
    `monitor_scoreboard_connection_TB4(2,1600,250);
    `monitor_scoreboard_connection_TB4(2,1601,251);
    `monitor_scoreboard_connection_TB4(2,1602,252);
    `monitor_scoreboard_connection_TB4(2,1603,253);
    `monitor_scoreboard_connection_TB4(2,1604,254);
    `monitor_scoreboard_connection_TB4(2,1605,255);
    `monitor_scoreboard_connection_TB4(2,1606,256);
    `monitor_scoreboard_connection_TB4(2,1607,257);
    `monitor_scoreboard_connection_TB4(2,1608,258);
    `monitor_scoreboard_connection_TB4(2,1609,259);
    `monitor_scoreboard_connection_TB4(2,1610,260);
    `monitor_scoreboard_connection_TB4(2,1611,261);
    `monitor_scoreboard_connection_TB4(2,1612,262);
    `monitor_scoreboard_connection_TB4(2,1613,263);
    `monitor_scoreboard_connection_TB4(2,1614,264);
    `monitor_scoreboard_connection_TB4(2,1615,265);
    `monitor_scoreboard_connection_TB4(2,1616,266);
    `monitor_scoreboard_connection_TB4(2,1617,267);
    `monitor_scoreboard_connection_TB4(2,1618,268);
    `monitor_scoreboard_connection_TB4(2,1619,269);
    `monitor_scoreboard_connection_TB4(2,1620,270);
    `monitor_scoreboard_connection_TB4(2,1621,271);
    `monitor_scoreboard_connection_TB4(2,1622,272);
    `monitor_scoreboard_connection_TB4(2,1623,273);
    `monitor_scoreboard_connection_TB4(2,1624,274);
    `monitor_scoreboard_connection_TB4(2,1625,275);
    `monitor_scoreboard_connection_TB4(2,1626,276);
    `monitor_scoreboard_connection_TB4(2,1627,277);
    `monitor_scoreboard_connection_TB4(2,1628,278);
    `monitor_scoreboard_connection_TB4(2,1629,279);
    `monitor_scoreboard_connection_TB4(2,1630,280);
    `monitor_scoreboard_connection_TB4(2,1631,281);
    `monitor_scoreboard_connection_TB4(2,1632,282);
    `monitor_scoreboard_connection_TB4(2,1633,283);
    `monitor_scoreboard_connection_TB4(2,1634,284);
    `monitor_scoreboard_connection_TB4(2,1635,285);
    `monitor_scoreboard_connection_TB4(2,1636,286);
    `monitor_scoreboard_connection_TB4(2,1637,287);
    `monitor_scoreboard_connection_TB4(2,1638,288);
    `monitor_scoreboard_connection_TB4(2,1639,289);
    `monitor_scoreboard_connection_TB4(2,1640,290);
    `monitor_scoreboard_connection_TB4(2,1641,291);
    `monitor_scoreboard_connection_TB4(2,1642,292);
    `monitor_scoreboard_connection_TB4(2,1643,293);
    `monitor_scoreboard_connection_TB4(2,1644,294);
    `monitor_scoreboard_connection_TB4(2,1645,295);
    `monitor_scoreboard_connection_TB4(2,1646,296);
    `monitor_scoreboard_connection_TB4(2,1647,297);
    `monitor_scoreboard_connection_TB4(2,1648,298);
    `monitor_scoreboard_connection_TB4(2,1649,299);
    `monitor_scoreboard_connection_TB4(2,1650,300);
    `monitor_scoreboard_connection_TB4(2,1651,301);
    `monitor_scoreboard_connection_TB4(2,1652,302);
    `monitor_scoreboard_connection_TB4(2,1653,303);
    `monitor_scoreboard_connection_TB4(2,1654,304);
    `monitor_scoreboard_connection_TB4(2,1655,305);
    `monitor_scoreboard_connection_TB4(2,1656,306);
    `monitor_scoreboard_connection_TB4(2,1657,307);
    `monitor_scoreboard_connection_TB4(2,1658,308);
    `monitor_scoreboard_connection_TB4(2,1659,309);
    `monitor_scoreboard_connection_TB4(2,1660,310);
    `monitor_scoreboard_connection_TB4(2,1661,311);
    `monitor_scoreboard_connection_TB4(2,1662,312);
    `monitor_scoreboard_connection_TB4(2,1663,313);
    `monitor_scoreboard_connection_TB4(2,1664,314);
    `monitor_scoreboard_connection_TB4(2,1665,315);
    `monitor_scoreboard_connection_TB4(2,1666,316);
    `monitor_scoreboard_connection_TB4(2,1667,317);
    `monitor_scoreboard_connection_TB4(2,1668,318);
    `monitor_scoreboard_connection_TB4(2,1669,319);
    `monitor_scoreboard_connection_TB4(2,1670,320);
    `monitor_scoreboard_connection_TB4(2,1671,321);
    `monitor_scoreboard_connection_TB4(2,1672,322);
    `monitor_scoreboard_connection_TB4(2,1673,323);
    `monitor_scoreboard_connection_TB4(2,1674,324);
    `monitor_scoreboard_connection_TB4(2,1675,325);
    `monitor_scoreboard_connection_TB4(2,1676,326);
    `monitor_scoreboard_connection_TB4(2,1677,327);
    `monitor_scoreboard_connection_TB4(2,1678,328);
    `monitor_scoreboard_connection_TB4(2,1679,329);
    `monitor_scoreboard_connection_TB4(2,1680,330);
    `monitor_scoreboard_connection_TB4(2,1681,331);
    `monitor_scoreboard_connection_TB4(2,1682,332);
    `monitor_scoreboard_connection_TB4(2,1683,333);
    `monitor_scoreboard_connection_TB4(2,1684,334);
    `monitor_scoreboard_connection_TB4(2,1685,335);
    `monitor_scoreboard_connection_TB4(2,1686,336);
    `monitor_scoreboard_connection_TB4(2,1687,337);
    `monitor_scoreboard_connection_TB4(2,1688,338);
    `monitor_scoreboard_connection_TB4(2,1689,339);
    `monitor_scoreboard_connection_TB4(2,1690,340);
    `monitor_scoreboard_connection_TB4(2,1691,341);
    `monitor_scoreboard_connection_TB4(2,1692,342);
    `monitor_scoreboard_connection_TB4(2,1693,343);
    `monitor_scoreboard_connection_TB4(2,1694,344);
    `monitor_scoreboard_connection_TB4(2,1695,345);
    `monitor_scoreboard_connection_TB4(2,1696,346);
    `monitor_scoreboard_connection_TB4(2,1697,347);
    `monitor_scoreboard_connection_TB4(2,1698,348);
    `monitor_scoreboard_connection_TB4(2,1699,349);
    `monitor_scoreboard_connection_TB4(2,1700,350);
    `monitor_scoreboard_connection_TB4(2,1701,351);
    `monitor_scoreboard_connection_TB4(2,1702,352);
    `monitor_scoreboard_connection_TB4(2,1703,353);
    `monitor_scoreboard_connection_TB4(2,1704,354);
    `monitor_scoreboard_connection_TB4(2,1705,355);
    `monitor_scoreboard_connection_TB4(2,1706,356);
    `monitor_scoreboard_connection_TB4(2,1707,357);
    `monitor_scoreboard_connection_TB4(2,1708,358);
    `monitor_scoreboard_connection_TB4(2,1709,359);
    `monitor_scoreboard_connection_TB4(2,1710,360);
    `monitor_scoreboard_connection_TB4(2,1711,361);
    `monitor_scoreboard_connection_TB4(2,1712,362);
    `monitor_scoreboard_connection_TB4(2,1713,363);
    `monitor_scoreboard_connection_TB4(2,1714,364);
    `monitor_scoreboard_connection_TB4(2,1715,365);
    `monitor_scoreboard_connection_TB4(2,1716,366);
    `monitor_scoreboard_connection_TB4(2,1717,367);
    `monitor_scoreboard_connection_TB4(2,1718,368);
    `monitor_scoreboard_connection_TB4(2,1719,369);
    `monitor_scoreboard_connection_TB4(2,1720,370);
    `monitor_scoreboard_connection_TB4(2,1721,371);
    `monitor_scoreboard_connection_TB4(2,1722,372);
    `monitor_scoreboard_connection_TB4(2,1723,373);
    `monitor_scoreboard_connection_TB4(2,1724,374);
    `monitor_scoreboard_connection_TB4(2,1725,375);
    `monitor_scoreboard_connection_TB4(2,1726,376);
    `monitor_scoreboard_connection_TB4(2,1727,377);
    `monitor_scoreboard_connection_TB4(2,1728,378);
    `monitor_scoreboard_connection_TB4(2,1729,379);
    `monitor_scoreboard_connection_TB4(2,1730,380);
    `monitor_scoreboard_connection_TB4(2,1731,381);
    `monitor_scoreboard_connection_TB4(2,1732,382);
    `monitor_scoreboard_connection_TB4(2,1733,383);
    `monitor_scoreboard_connection_TB4(2,1734,384);
    `monitor_scoreboard_connection_TB4(2,1735,385);
    `monitor_scoreboard_connection_TB4(2,1736,386);
    `monitor_scoreboard_connection_TB4(2,1737,387);
    `monitor_scoreboard_connection_TB4(2,1738,388);
    `monitor_scoreboard_connection_TB4(2,1739,389);
    `monitor_scoreboard_connection_TB4(2,1740,390);
    `monitor_scoreboard_connection_TB4(2,1741,391);
    `monitor_scoreboard_connection_TB4(2,1742,392);
    `monitor_scoreboard_connection_TB4(2,1743,393);
    `monitor_scoreboard_connection_TB4(2,1744,394);
    `monitor_scoreboard_connection_TB4(2,1745,395);
    `monitor_scoreboard_connection_TB4(2,1746,396);
    `monitor_scoreboard_connection_TB4(2,1747,397);
    `monitor_scoreboard_connection_TB4(2,1748,398);
    `monitor_scoreboard_connection_TB4(2,1749,399);
    `monitor_scoreboard_connection_TB4(2,1750,400);
    `monitor_scoreboard_connection_TB4(2,1751,401);
    `monitor_scoreboard_connection_TB4(2,1752,402);
    `monitor_scoreboard_connection_TB4(2,1753,403);
    `monitor_scoreboard_connection_TB4(2,1754,404);
    `monitor_scoreboard_connection_TB4(2,1755,405);
    `monitor_scoreboard_connection_TB4(2,1756,406);
    `monitor_scoreboard_connection_TB4(2,1757,407);
    `monitor_scoreboard_connection_TB4(2,1758,408);
    `monitor_scoreboard_connection_TB4(2,1759,409);
    `monitor_scoreboard_connection_TB4(2,1760,410);
    `monitor_scoreboard_connection_TB4(2,1761,411);
    `monitor_scoreboard_connection_TB4(2,1762,412);
    `monitor_scoreboard_connection_TB4(2,1763,413);
    `monitor_scoreboard_connection_TB4(2,1764,414);
    `monitor_scoreboard_connection_TB4(2,1765,415);
    `monitor_scoreboard_connection_TB4(2,1766,416);
    `monitor_scoreboard_connection_TB4(2,1767,417);
    `monitor_scoreboard_connection_TB4(2,1768,418);
    `monitor_scoreboard_connection_TB4(2,1769,419);
    `monitor_scoreboard_connection_TB4(2,1770,420);
    `monitor_scoreboard_connection_TB4(2,1771,421);
    `monitor_scoreboard_connection_TB4(2,1772,422);
    `monitor_scoreboard_connection_TB4(2,1773,423);
    `monitor_scoreboard_connection_TB4(2,1774,424);
    `monitor_scoreboard_connection_TB4(2,1775,425);
    `monitor_scoreboard_connection_TB4(2,1776,426);
    `monitor_scoreboard_connection_TB4(2,1777,427);
    `monitor_scoreboard_connection_TB4(2,1778,428);
    `monitor_scoreboard_connection_TB4(2,1779,429);
    `monitor_scoreboard_connection_TB4(2,1780,430);
    `monitor_scoreboard_connection_TB4(2,1781,431);
    `monitor_scoreboard_connection_TB4(2,1782,432);
    `monitor_scoreboard_connection_TB4(2,1783,433);
    `monitor_scoreboard_connection_TB4(2,1784,434);
    `monitor_scoreboard_connection_TB4(2,1785,435);
    `monitor_scoreboard_connection_TB4(2,1786,436);
    `monitor_scoreboard_connection_TB4(2,1787,437);
    `monitor_scoreboard_connection_TB4(2,1788,438);
    `monitor_scoreboard_connection_TB4(2,1789,439);
    `monitor_scoreboard_connection_TB4(2,1790,440);
    `monitor_scoreboard_connection_TB4(2,1791,441);
    `monitor_scoreboard_connection_TB4(2,1792,442);
    `monitor_scoreboard_connection_TB4(2,1793,443);
    `monitor_scoreboard_connection_TB4(2,1794,444);
    `monitor_scoreboard_connection_TB4(2,1795,445);
    `monitor_scoreboard_connection_TB4(2,1796,446);
    `monitor_scoreboard_connection_TB4(2,1797,447);
    `monitor_scoreboard_connection_TB4(2,1798,448);
    `monitor_scoreboard_connection_TB4(2,1799,449);
    `monitor_scoreboard_connection_TB4(3,1800,0);
    `monitor_scoreboard_connection_TB4(3,1801,1);
    `monitor_scoreboard_connection_TB4(3,1802,2);
    `monitor_scoreboard_connection_TB4(3,1803,3);
    `monitor_scoreboard_connection_TB4(3,1804,4);
    `monitor_scoreboard_connection_TB4(3,1805,5);
    `monitor_scoreboard_connection_TB4(3,1806,6);
    `monitor_scoreboard_connection_TB4(3,1807,7);
    `monitor_scoreboard_connection_TB4(3,1808,8);
    `monitor_scoreboard_connection_TB4(3,1809,9);
    `monitor_scoreboard_connection_TB4(3,1810,10);
    `monitor_scoreboard_connection_TB4(3,1811,11);
    `monitor_scoreboard_connection_TB4(3,1812,12);
    `monitor_scoreboard_connection_TB4(3,1813,13);
    `monitor_scoreboard_connection_TB4(3,1814,14);
    `monitor_scoreboard_connection_TB4(3,1815,15);
    `monitor_scoreboard_connection_TB4(3,1816,16);
    `monitor_scoreboard_connection_TB4(3,1817,17);
    `monitor_scoreboard_connection_TB4(3,1818,18);
    `monitor_scoreboard_connection_TB4(3,1819,19);
    `monitor_scoreboard_connection_TB4(3,1820,20);
    `monitor_scoreboard_connection_TB4(3,1821,21);
    `monitor_scoreboard_connection_TB4(3,1822,22);
    `monitor_scoreboard_connection_TB4(3,1823,23);
    `monitor_scoreboard_connection_TB4(3,1824,24);
    `monitor_scoreboard_connection_TB4(3,1825,25);
    `monitor_scoreboard_connection_TB4(3,1826,26);
    `monitor_scoreboard_connection_TB4(3,1827,27);
    `monitor_scoreboard_connection_TB4(3,1828,28);
    `monitor_scoreboard_connection_TB4(3,1829,29);
    `monitor_scoreboard_connection_TB4(3,1830,30);
    `monitor_scoreboard_connection_TB4(3,1831,31);
    `monitor_scoreboard_connection_TB4(3,1832,32);
    `monitor_scoreboard_connection_TB4(3,1833,33);
    `monitor_scoreboard_connection_TB4(3,1834,34);
    `monitor_scoreboard_connection_TB4(3,1835,35);
    `monitor_scoreboard_connection_TB4(3,1836,36);
    `monitor_scoreboard_connection_TB4(3,1837,37);
    `monitor_scoreboard_connection_TB4(3,1838,38);
    `monitor_scoreboard_connection_TB4(3,1839,39);
    `monitor_scoreboard_connection_TB4(3,1840,40);
    `monitor_scoreboard_connection_TB4(3,1841,41);
    `monitor_scoreboard_connection_TB4(3,1842,42);
    `monitor_scoreboard_connection_TB4(3,1843,43);
    `monitor_scoreboard_connection_TB4(3,1844,44);
    `monitor_scoreboard_connection_TB4(3,1845,45);
    `monitor_scoreboard_connection_TB4(3,1846,46);
    `monitor_scoreboard_connection_TB4(3,1847,47);
    `monitor_scoreboard_connection_TB4(3,1848,48);
    `monitor_scoreboard_connection_TB4(3,1849,49);
    `monitor_scoreboard_connection_TB4(3,1850,50);
    `monitor_scoreboard_connection_TB4(3,1851,51);
    `monitor_scoreboard_connection_TB4(3,1852,52);
    `monitor_scoreboard_connection_TB4(3,1853,53);
    `monitor_scoreboard_connection_TB4(3,1854,54);
    `monitor_scoreboard_connection_TB4(3,1855,55);
    `monitor_scoreboard_connection_TB4(3,1856,56);
    `monitor_scoreboard_connection_TB4(3,1857,57);
    `monitor_scoreboard_connection_TB4(3,1858,58);
    `monitor_scoreboard_connection_TB4(3,1859,59);
    `monitor_scoreboard_connection_TB4(3,1860,60);
    `monitor_scoreboard_connection_TB4(3,1861,61);
    `monitor_scoreboard_connection_TB4(3,1862,62);
    `monitor_scoreboard_connection_TB4(3,1863,63);
    `monitor_scoreboard_connection_TB4(3,1864,64);
    `monitor_scoreboard_connection_TB4(3,1865,65);
    `monitor_scoreboard_connection_TB4(3,1866,66);
    `monitor_scoreboard_connection_TB4(3,1867,67);
    `monitor_scoreboard_connection_TB4(3,1868,68);
    `monitor_scoreboard_connection_TB4(3,1869,69);
    `monitor_scoreboard_connection_TB4(3,1870,70);
    `monitor_scoreboard_connection_TB4(3,1871,71);
    `monitor_scoreboard_connection_TB4(3,1872,72);
    `monitor_scoreboard_connection_TB4(3,1873,73);
    `monitor_scoreboard_connection_TB4(3,1874,74);
    `monitor_scoreboard_connection_TB4(3,1875,75);
    `monitor_scoreboard_connection_TB4(3,1876,76);
    `monitor_scoreboard_connection_TB4(3,1877,77);
    `monitor_scoreboard_connection_TB4(3,1878,78);
    `monitor_scoreboard_connection_TB4(3,1879,79);
    `monitor_scoreboard_connection_TB4(3,1880,80);
    `monitor_scoreboard_connection_TB4(3,1881,81);
    `monitor_scoreboard_connection_TB4(3,1882,82);
    `monitor_scoreboard_connection_TB4(3,1883,83);
    `monitor_scoreboard_connection_TB4(3,1884,84);
    `monitor_scoreboard_connection_TB4(3,1885,85);
    `monitor_scoreboard_connection_TB4(3,1886,86);
    `monitor_scoreboard_connection_TB4(3,1887,87);
    `monitor_scoreboard_connection_TB4(3,1888,88);
    `monitor_scoreboard_connection_TB4(3,1889,89);
    `monitor_scoreboard_connection_TB4(3,1890,90);
    `monitor_scoreboard_connection_TB4(3,1891,91);
    `monitor_scoreboard_connection_TB4(3,1892,92);
    `monitor_scoreboard_connection_TB4(3,1893,93);
    `monitor_scoreboard_connection_TB4(3,1894,94);
    `monitor_scoreboard_connection_TB4(3,1895,95);
    `monitor_scoreboard_connection_TB4(3,1896,96);
    `monitor_scoreboard_connection_TB4(3,1897,97);
    `monitor_scoreboard_connection_TB4(3,1898,98);
    `monitor_scoreboard_connection_TB4(3,1899,99);
    `monitor_scoreboard_connection_TB4(3,1900,100);
    `monitor_scoreboard_connection_TB4(3,1901,101);
    `monitor_scoreboard_connection_TB4(3,1902,102);
    `monitor_scoreboard_connection_TB4(3,1903,103);
    `monitor_scoreboard_connection_TB4(3,1904,104);
    `monitor_scoreboard_connection_TB4(3,1905,105);
    `monitor_scoreboard_connection_TB4(3,1906,106);
    `monitor_scoreboard_connection_TB4(3,1907,107);
    `monitor_scoreboard_connection_TB4(3,1908,108);
    `monitor_scoreboard_connection_TB4(3,1909,109);
    `monitor_scoreboard_connection_TB4(3,1910,110);
    `monitor_scoreboard_connection_TB4(3,1911,111);
    `monitor_scoreboard_connection_TB4(3,1912,112);
    `monitor_scoreboard_connection_TB4(3,1913,113);
    `monitor_scoreboard_connection_TB4(3,1914,114);
    `monitor_scoreboard_connection_TB4(3,1915,115);
    `monitor_scoreboard_connection_TB4(3,1916,116);
    `monitor_scoreboard_connection_TB4(3,1917,117);
    `monitor_scoreboard_connection_TB4(3,1918,118);
    `monitor_scoreboard_connection_TB4(3,1919,119);
    `monitor_scoreboard_connection_TB4(3,1920,120);
    `monitor_scoreboard_connection_TB4(3,1921,121);
    `monitor_scoreboard_connection_TB4(3,1922,122);
    `monitor_scoreboard_connection_TB4(3,1923,123);
    `monitor_scoreboard_connection_TB4(3,1924,124);
    `monitor_scoreboard_connection_TB4(3,1925,125);
    `monitor_scoreboard_connection_TB4(3,1926,126);
    `monitor_scoreboard_connection_TB4(3,1927,127);
    `monitor_scoreboard_connection_TB4(3,1928,128);
    `monitor_scoreboard_connection_TB4(3,1929,129);
    `monitor_scoreboard_connection_TB4(3,1930,130);
    `monitor_scoreboard_connection_TB4(3,1931,131);
    `monitor_scoreboard_connection_TB4(3,1932,132);
    `monitor_scoreboard_connection_TB4(3,1933,133);
    `monitor_scoreboard_connection_TB4(3,1934,134);
    `monitor_scoreboard_connection_TB4(3,1935,135);
    `monitor_scoreboard_connection_TB4(3,1936,136);
    `monitor_scoreboard_connection_TB4(3,1937,137);
    `monitor_scoreboard_connection_TB4(3,1938,138);
    `monitor_scoreboard_connection_TB4(3,1939,139);
    `monitor_scoreboard_connection_TB4(3,1940,140);
    `monitor_scoreboard_connection_TB4(3,1941,141);
    `monitor_scoreboard_connection_TB4(3,1942,142);
    `monitor_scoreboard_connection_TB4(3,1943,143);
    `monitor_scoreboard_connection_TB4(3,1944,144);
    `monitor_scoreboard_connection_TB4(3,1945,145);
    `monitor_scoreboard_connection_TB4(3,1946,146);
    `monitor_scoreboard_connection_TB4(3,1947,147);
    `monitor_scoreboard_connection_TB4(3,1948,148);
    `monitor_scoreboard_connection_TB4(3,1949,149);
    `monitor_scoreboard_connection_TB4(3,1950,150);
    `monitor_scoreboard_connection_TB4(3,1951,151);
    `monitor_scoreboard_connection_TB4(3,1952,152);
    `monitor_scoreboard_connection_TB4(3,1953,153);
    `monitor_scoreboard_connection_TB4(3,1954,154);
    `monitor_scoreboard_connection_TB4(3,1955,155);
    `monitor_scoreboard_connection_TB4(3,1956,156);
    `monitor_scoreboard_connection_TB4(3,1957,157);
    `monitor_scoreboard_connection_TB4(3,1958,158);
    `monitor_scoreboard_connection_TB4(3,1959,159);
    `monitor_scoreboard_connection_TB4(3,1960,160);
    `monitor_scoreboard_connection_TB4(3,1961,161);
    `monitor_scoreboard_connection_TB4(3,1962,162);
    `monitor_scoreboard_connection_TB4(3,1963,163);
    `monitor_scoreboard_connection_TB4(3,1964,164);
    `monitor_scoreboard_connection_TB4(3,1965,165);
    `monitor_scoreboard_connection_TB4(3,1966,166);
    `monitor_scoreboard_connection_TB4(3,1967,167);
    `monitor_scoreboard_connection_TB4(3,1968,168);
    `monitor_scoreboard_connection_TB4(3,1969,169);
    `monitor_scoreboard_connection_TB4(3,1970,170);
    `monitor_scoreboard_connection_TB4(3,1971,171);
    `monitor_scoreboard_connection_TB4(3,1972,172);
    `monitor_scoreboard_connection_TB4(3,1973,173);
    `monitor_scoreboard_connection_TB4(3,1974,174);
    `monitor_scoreboard_connection_TB4(3,1975,175);
    `monitor_scoreboard_connection_TB4(3,1976,176);
    `monitor_scoreboard_connection_TB4(3,1977,177);
    `monitor_scoreboard_connection_TB4(3,1978,178);
    `monitor_scoreboard_connection_TB4(3,1979,179);
    `monitor_scoreboard_connection_TB4(3,1980,180);
    `monitor_scoreboard_connection_TB4(3,1981,181);
    `monitor_scoreboard_connection_TB4(3,1982,182);
    `monitor_scoreboard_connection_TB4(3,1983,183);
    `monitor_scoreboard_connection_TB4(3,1984,184);
    `monitor_scoreboard_connection_TB4(3,1985,185);
    `monitor_scoreboard_connection_TB4(3,1986,186);
    `monitor_scoreboard_connection_TB4(3,1987,187);
    `monitor_scoreboard_connection_TB4(3,1988,188);
    `monitor_scoreboard_connection_TB4(3,1989,189);
    `monitor_scoreboard_connection_TB4(3,1990,190);
    `monitor_scoreboard_connection_TB4(3,1991,191);
    `monitor_scoreboard_connection_TB4(3,1992,192);
    `monitor_scoreboard_connection_TB4(3,1993,193);
    `monitor_scoreboard_connection_TB4(3,1994,194);
    `monitor_scoreboard_connection_TB4(3,1995,195);
    `monitor_scoreboard_connection_TB4(3,1996,196);
    `monitor_scoreboard_connection_TB4(3,1997,197);
    `monitor_scoreboard_connection_TB4(3,1998,198);
    `monitor_scoreboard_connection_TB4(3,1999,199);
    `monitor_scoreboard_connection_TB4(3,2000,200);
    `monitor_scoreboard_connection_TB4(3,2001,201);
    `monitor_scoreboard_connection_TB4(3,2002,202);
    `monitor_scoreboard_connection_TB4(3,2003,203);
    `monitor_scoreboard_connection_TB4(3,2004,204);
    `monitor_scoreboard_connection_TB4(3,2005,205);
    `monitor_scoreboard_connection_TB4(3,2006,206);
    `monitor_scoreboard_connection_TB4(3,2007,207);
    `monitor_scoreboard_connection_TB4(3,2008,208);
    `monitor_scoreboard_connection_TB4(3,2009,209);
    `monitor_scoreboard_connection_TB4(3,2010,210);
    `monitor_scoreboard_connection_TB4(3,2011,211);
    `monitor_scoreboard_connection_TB4(3,2012,212);
    `monitor_scoreboard_connection_TB4(3,2013,213);
    `monitor_scoreboard_connection_TB4(3,2014,214);
    `monitor_scoreboard_connection_TB4(3,2015,215);
    `monitor_scoreboard_connection_TB4(3,2016,216);
    `monitor_scoreboard_connection_TB4(3,2017,217);
    `monitor_scoreboard_connection_TB4(3,2018,218);
    `monitor_scoreboard_connection_TB4(3,2019,219);
    `monitor_scoreboard_connection_TB4(3,2020,220);
    `monitor_scoreboard_connection_TB4(3,2021,221);
    `monitor_scoreboard_connection_TB4(3,2022,222);
    `monitor_scoreboard_connection_TB4(3,2023,223);
    `monitor_scoreboard_connection_TB4(3,2024,224);
    `monitor_scoreboard_connection_TB4(3,2025,225);
    `monitor_scoreboard_connection_TB4(3,2026,226);
    `monitor_scoreboard_connection_TB4(3,2027,227);
    `monitor_scoreboard_connection_TB4(3,2028,228);
    `monitor_scoreboard_connection_TB4(3,2029,229);
    `monitor_scoreboard_connection_TB4(3,2030,230);
    `monitor_scoreboard_connection_TB4(3,2031,231);
    `monitor_scoreboard_connection_TB4(3,2032,232);
    `monitor_scoreboard_connection_TB4(3,2033,233);
    `monitor_scoreboard_connection_TB4(3,2034,234);
    `monitor_scoreboard_connection_TB4(3,2035,235);
    `monitor_scoreboard_connection_TB4(3,2036,236);
    `monitor_scoreboard_connection_TB4(3,2037,237);
    `monitor_scoreboard_connection_TB4(3,2038,238);
    `monitor_scoreboard_connection_TB4(3,2039,239);
    `monitor_scoreboard_connection_TB4(3,2040,240);
    `monitor_scoreboard_connection_TB4(3,2041,241);
    `monitor_scoreboard_connection_TB4(3,2042,242);
    `monitor_scoreboard_connection_TB4(3,2043,243);
    `monitor_scoreboard_connection_TB4(3,2044,244);
    `monitor_scoreboard_connection_TB4(3,2045,245);
    `monitor_scoreboard_connection_TB4(3,2046,246);
    `monitor_scoreboard_connection_TB4(3,2047,247);
    `monitor_scoreboard_upstream_connection(16);
    `monitor_scoreboard_upstream_connection(17);
    `monitor_scoreboard_upstream_connection(18);
    `monitor_scoreboard_upstream_connection(19);
    `monitor_scoreboard_upstream_connection(20);
    `monitor_scoreboard_upstream_connection(21);
    `monitor_scoreboard_upstream_connection(22);
    `monitor_scoreboard_upstream_connection(23);
    `monitor_scoreboard_upstream_connection(24);
    `monitor_scoreboard_upstream_connection(25);
    `monitor_scoreboard_upstream_connection(26);
    `monitor_scoreboard_upstream_connection(27);
    `monitor_scoreboard_upstream_connection(28);
    `monitor_scoreboard_upstream_connection(29);
    `monitor_scoreboard_upstream_connection(30);
    `monitor_scoreboard_upstream_connection(31);
    `monitor_scoreboard_upstream_connection(32);
    `monitor_scoreboard_upstream_connection(33);
    `monitor_scoreboard_upstream_connection(34);
    `monitor_scoreboard_upstream_connection(35);
    `monitor_scoreboard_upstream_connection(36);
    `monitor_scoreboard_upstream_connection(37);
    `monitor_scoreboard_upstream_connection(38);
    `monitor_scoreboard_upstream_connection(39);
    `monitor_scoreboard_upstream_connection(40);
    `monitor_scoreboard_upstream_connection(41);
    `monitor_scoreboard_upstream_connection(42);
    `monitor_scoreboard_upstream_connection(43);
    `monitor_scoreboard_upstream_connection(44);
    `monitor_scoreboard_upstream_connection(45);
    `monitor_scoreboard_upstream_connection(46);
    `monitor_scoreboard_upstream_connection(47);
    `monitor_scoreboard_upstream_connection(48);
    `monitor_scoreboard_upstream_connection(49);
    `monitor_scoreboard_upstream_connection(50);
    `monitor_scoreboard_upstream_connection(51);
    `monitor_scoreboard_upstream_connection(52);
    `monitor_scoreboard_upstream_connection(53);
    `monitor_scoreboard_upstream_connection(54);
    `monitor_scoreboard_upstream_connection(55);
    `monitor_scoreboard_upstream_connection(56);
    `monitor_scoreboard_upstream_connection(57);
    `monitor_scoreboard_upstream_connection(58);
    `monitor_scoreboard_upstream_connection(59);
    `monitor_scoreboard_upstream_connection(60);
    `monitor_scoreboard_upstream_connection(61);
    `monitor_scoreboard_upstream_connection(62);
    `monitor_scoreboard_upstream_connection(63);
    `monitor_scoreboard_upstream_connection(64);
    `monitor_scoreboard_upstream_connection(65);
    `monitor_scoreboard_upstream_connection(66);
    `monitor_scoreboard_upstream_connection(67);
    `monitor_scoreboard_upstream_connection(68);
    `monitor_scoreboard_upstream_connection(69);
    `monitor_scoreboard_upstream_connection(70);
    `monitor_scoreboard_upstream_connection(71);
    `monitor_scoreboard_upstream_connection(72);
    `monitor_scoreboard_upstream_connection(73);
    `monitor_scoreboard_upstream_connection(74);
    `monitor_scoreboard_upstream_connection(75);
    `monitor_scoreboard_upstream_connection(76);
    `monitor_scoreboard_upstream_connection(77);
    `monitor_scoreboard_upstream_connection(78);
    `monitor_scoreboard_upstream_connection(79);
    `monitor_scoreboard_upstream_connection(80);
    `monitor_scoreboard_upstream_connection(81);
    `monitor_scoreboard_upstream_connection(82);
    `monitor_scoreboard_upstream_connection(83);
    `monitor_scoreboard_upstream_connection(84);
    `monitor_scoreboard_upstream_connection(85);
    `monitor_scoreboard_upstream_connection(86);
    `monitor_scoreboard_upstream_connection(87);
    `monitor_scoreboard_upstream_connection(88);
    `monitor_scoreboard_upstream_connection(89);
    `monitor_scoreboard_upstream_connection(90);
    `monitor_scoreboard_upstream_connection(91);
    `monitor_scoreboard_upstream_connection(92);
    `monitor_scoreboard_upstream_connection(93);
    `monitor_scoreboard_upstream_connection(94);
    `monitor_scoreboard_upstream_connection(95);
    `monitor_scoreboard_upstream_connection(96);
    `monitor_scoreboard_upstream_connection(97);
    `monitor_scoreboard_upstream_connection(98);
    `monitor_scoreboard_upstream_connection(99);
    `monitor_scoreboard_upstream_connection(100);
    `monitor_scoreboard_upstream_connection(101);
    `monitor_scoreboard_upstream_connection(102);
    `monitor_scoreboard_upstream_connection(103);
    `monitor_scoreboard_upstream_connection(104);
    `monitor_scoreboard_upstream_connection(105);
    `monitor_scoreboard_upstream_connection(106);
    `monitor_scoreboard_upstream_connection(107);
    `monitor_scoreboard_upstream_connection(108);
    `monitor_scoreboard_upstream_connection(109);
    `monitor_scoreboard_upstream_connection(110);
    `monitor_scoreboard_upstream_connection(111);
    `monitor_scoreboard_upstream_connection(112);
    `monitor_scoreboard_upstream_connection(113);
    `monitor_scoreboard_upstream_connection(114);
    `monitor_scoreboard_upstream_connection(115);
    `monitor_scoreboard_upstream_connection(116);
    `monitor_scoreboard_upstream_connection(117);
    `monitor_scoreboard_upstream_connection(118);
    `monitor_scoreboard_upstream_connection(119);
    `monitor_scoreboard_upstream_connection(120);
    `monitor_scoreboard_upstream_connection(121);
    `monitor_scoreboard_upstream_connection(122);
    `monitor_scoreboard_upstream_connection(123);
    `monitor_scoreboard_upstream_connection(124);
    `monitor_scoreboard_upstream_connection(125);
    `monitor_scoreboard_upstream_connection(126);
    `monitor_scoreboard_upstream_connection(127);
    `monitor_scoreboard_upstream_connection(128);
    `monitor_scoreboard_upstream_connection(129);
    `monitor_scoreboard_upstream_connection(130);
    `monitor_scoreboard_upstream_connection(131);
    `monitor_scoreboard_upstream_connection(132);
    `monitor_scoreboard_upstream_connection(133);
    `monitor_scoreboard_upstream_connection(134);
    `monitor_scoreboard_upstream_connection(135);
    `monitor_scoreboard_upstream_connection(136);
    `monitor_scoreboard_upstream_connection(137);
    `monitor_scoreboard_upstream_connection(138);
    `monitor_scoreboard_upstream_connection(139);
    `monitor_scoreboard_upstream_connection(140);
    `monitor_scoreboard_upstream_connection(141);
    `monitor_scoreboard_upstream_connection(142);
    `monitor_scoreboard_upstream_connection(143);
    `monitor_scoreboard_upstream_connection(144);
    `monitor_scoreboard_upstream_connection(145);
    `monitor_scoreboard_upstream_connection(146);
    `monitor_scoreboard_upstream_connection(147);
    `monitor_scoreboard_upstream_connection(148);
    `monitor_scoreboard_upstream_connection(149);
    `monitor_scoreboard_upstream_connection(150);
    `monitor_scoreboard_upstream_connection(151);
    `monitor_scoreboard_upstream_connection(152);
    `monitor_scoreboard_upstream_connection(153);
    `monitor_scoreboard_upstream_connection(154);
    `monitor_scoreboard_upstream_connection(155);
    `monitor_scoreboard_upstream_connection(156);
    `monitor_scoreboard_upstream_connection(157);
    `monitor_scoreboard_upstream_connection(158);
    `monitor_scoreboard_upstream_connection(159);
    `monitor_scoreboard_upstream_connection(160);
    `monitor_scoreboard_upstream_connection(161);
    `monitor_scoreboard_upstream_connection(162);
    `monitor_scoreboard_upstream_connection(163);
    `monitor_scoreboard_upstream_connection(164);
    `monitor_scoreboard_upstream_connection(165);
    `monitor_scoreboard_upstream_connection(166);
    `monitor_scoreboard_upstream_connection(167);
    `monitor_scoreboard_upstream_connection(168);
    `monitor_scoreboard_upstream_connection(169);
    `monitor_scoreboard_upstream_connection(170);
    `monitor_scoreboard_upstream_connection(171);
    `monitor_scoreboard_upstream_connection(172);
    `monitor_scoreboard_upstream_connection(173);
    `monitor_scoreboard_upstream_connection(174);
    `monitor_scoreboard_upstream_connection(175);
    `monitor_scoreboard_upstream_connection(176);
    `monitor_scoreboard_upstream_connection(177);
    `monitor_scoreboard_upstream_connection(178);
    `monitor_scoreboard_upstream_connection(179);
    `monitor_scoreboard_upstream_connection(180);
    `monitor_scoreboard_upstream_connection(181);
    `monitor_scoreboard_upstream_connection(182);
    `monitor_scoreboard_upstream_connection(183);
    `monitor_scoreboard_upstream_connection(184);
    `monitor_scoreboard_upstream_connection(185);
    `monitor_scoreboard_upstream_connection(186);
    `monitor_scoreboard_upstream_connection(187);
    `monitor_scoreboard_upstream_connection(188);
    `monitor_scoreboard_upstream_connection(189);
    `monitor_scoreboard_upstream_connection(190);
    `monitor_scoreboard_upstream_connection(191);
    `monitor_scoreboard_upstream_connection(192);
    `monitor_scoreboard_upstream_connection(193);
    `monitor_scoreboard_upstream_connection(194);
    `monitor_scoreboard_upstream_connection(195);
    `monitor_scoreboard_upstream_connection(196);
    `monitor_scoreboard_upstream_connection(197);
    `monitor_scoreboard_upstream_connection(198);
    `monitor_scoreboard_upstream_connection(199);
    `monitor_scoreboard_upstream_connection(200);
    `monitor_scoreboard_upstream_connection(201);
    `monitor_scoreboard_upstream_connection(202);
    `monitor_scoreboard_upstream_connection(203);
    `monitor_scoreboard_upstream_connection(204);
    `monitor_scoreboard_upstream_connection(205);
    `monitor_scoreboard_upstream_connection(206);
    `monitor_scoreboard_upstream_connection(207);
    `monitor_scoreboard_upstream_connection(208);
    `monitor_scoreboard_upstream_connection(209);
    `monitor_scoreboard_upstream_connection(210);
    `monitor_scoreboard_upstream_connection(211);
    `monitor_scoreboard_upstream_connection(212);
    `monitor_scoreboard_upstream_connection(213);
    `monitor_scoreboard_upstream_connection(214);
    `monitor_scoreboard_upstream_connection(215);
    `monitor_scoreboard_upstream_connection(216);
    `monitor_scoreboard_upstream_connection(217);
    `monitor_scoreboard_upstream_connection(218);
    `monitor_scoreboard_upstream_connection(219);
    `monitor_scoreboard_upstream_connection(220);
    `monitor_scoreboard_upstream_connection(221);
    `monitor_scoreboard_upstream_connection(222);
    `monitor_scoreboard_upstream_connection(223);
    `monitor_scoreboard_upstream_connection(224);
    `monitor_scoreboard_upstream_connection(225);
    `monitor_scoreboard_upstream_connection(226);
    `monitor_scoreboard_upstream_connection(227);
    `monitor_scoreboard_upstream_connection(228);
    `monitor_scoreboard_upstream_connection(229);
    `monitor_scoreboard_upstream_connection(230);
    `monitor_scoreboard_upstream_connection(231);
    `monitor_scoreboard_upstream_connection(232);
    `monitor_scoreboard_upstream_connection(233);
    `monitor_scoreboard_upstream_connection(234);
    `monitor_scoreboard_upstream_connection(235);
    `monitor_scoreboard_upstream_connection(236);
    `monitor_scoreboard_upstream_connection(237);
    `monitor_scoreboard_upstream_connection(238);
    `monitor_scoreboard_upstream_connection(239);
    `monitor_scoreboard_upstream_connection(240);
    `monitor_scoreboard_upstream_connection(241);
    `monitor_scoreboard_upstream_connection(242);
    `monitor_scoreboard_upstream_connection(243);
    `monitor_scoreboard_upstream_connection(244);
    `monitor_scoreboard_upstream_connection(245);
    `monitor_scoreboard_upstream_connection(246);
    `monitor_scoreboard_upstream_connection(247);
    `monitor_scoreboard_upstream_connection(248);
    `monitor_scoreboard_upstream_connection(249);
    `monitor_scoreboard_upstream_connection(250);
    `monitor_scoreboard_upstream_connection(251);
    `monitor_scoreboard_upstream_connection(252);
    `monitor_scoreboard_upstream_connection(253);
    `monitor_scoreboard_upstream_connection(254);
    `monitor_scoreboard_upstream_connection(255);
    `monitor_scoreboard_upstream_connection(256);
    `monitor_scoreboard_upstream_connection(257);
    `monitor_scoreboard_upstream_connection(258);
    `monitor_scoreboard_upstream_connection(259);
    `monitor_scoreboard_upstream_connection(260);
    `monitor_scoreboard_upstream_connection(261);
    `monitor_scoreboard_upstream_connection(262);
    `monitor_scoreboard_upstream_connection(263);
    `monitor_scoreboard_upstream_connection(264);
    `monitor_scoreboard_upstream_connection(265);
    `monitor_scoreboard_upstream_connection(266);
    `monitor_scoreboard_upstream_connection(267);
    `monitor_scoreboard_upstream_connection(268);
    `monitor_scoreboard_upstream_connection(269);
    `monitor_scoreboard_upstream_connection(270);
    `monitor_scoreboard_upstream_connection(271);
    `monitor_scoreboard_upstream_connection(272);
    `monitor_scoreboard_upstream_connection(273);
    `monitor_scoreboard_upstream_connection(274);
    `monitor_scoreboard_upstream_connection(275);
    `monitor_scoreboard_upstream_connection(276);
    `monitor_scoreboard_upstream_connection(277);
    `monitor_scoreboard_upstream_connection(278);
    `monitor_scoreboard_upstream_connection(279);
    `monitor_scoreboard_upstream_connection(280);
    `monitor_scoreboard_upstream_connection(281);
    `monitor_scoreboard_upstream_connection(282);
    `monitor_scoreboard_upstream_connection(283);
    `monitor_scoreboard_upstream_connection(284);
    `monitor_scoreboard_upstream_connection(285);
    `monitor_scoreboard_upstream_connection(286);
    `monitor_scoreboard_upstream_connection(287);
    `monitor_scoreboard_upstream_connection(288);
    `monitor_scoreboard_upstream_connection(289);
    `monitor_scoreboard_upstream_connection(290);
    `monitor_scoreboard_upstream_connection(291);
    `monitor_scoreboard_upstream_connection(292);
    `monitor_scoreboard_upstream_connection(293);
    `monitor_scoreboard_upstream_connection(294);
    `monitor_scoreboard_upstream_connection(295);
    `monitor_scoreboard_upstream_connection(296);
    `monitor_scoreboard_upstream_connection(297);
    `monitor_scoreboard_upstream_connection(298);
    `monitor_scoreboard_upstream_connection(299);
    `monitor_scoreboard_upstream_connection(300);
    `monitor_scoreboard_upstream_connection(301);
    `monitor_scoreboard_upstream_connection(302);
    `monitor_scoreboard_upstream_connection(303);
    `monitor_scoreboard_upstream_connection(304);
    `monitor_scoreboard_upstream_connection(305);
    `monitor_scoreboard_upstream_connection(306);
    `monitor_scoreboard_upstream_connection(307);
    `monitor_scoreboard_upstream_connection(308);
    `monitor_scoreboard_upstream_connection(309);
    `monitor_scoreboard_upstream_connection(310);
    `monitor_scoreboard_upstream_connection(311);
    `monitor_scoreboard_upstream_connection(312);
    `monitor_scoreboard_upstream_connection(313);
    `monitor_scoreboard_upstream_connection(314);
    `monitor_scoreboard_upstream_connection(315);
    `monitor_scoreboard_upstream_connection(316);
    `monitor_scoreboard_upstream_connection(317);
    `monitor_scoreboard_upstream_connection(318);
    `monitor_scoreboard_upstream_connection(319);
    `monitor_scoreboard_upstream_connection(320);
    `monitor_scoreboard_upstream_connection(321);
    `monitor_scoreboard_upstream_connection(322);
    `monitor_scoreboard_upstream_connection(323);
    `monitor_scoreboard_upstream_connection(324);
    `monitor_scoreboard_upstream_connection(325);
    `monitor_scoreboard_upstream_connection(326);
    `monitor_scoreboard_upstream_connection(327);
    `monitor_scoreboard_upstream_connection(328);
    `monitor_scoreboard_upstream_connection(329);
    `monitor_scoreboard_upstream_connection(330);
    `monitor_scoreboard_upstream_connection(331);
    `monitor_scoreboard_upstream_connection(332);
    `monitor_scoreboard_upstream_connection(333);
    `monitor_scoreboard_upstream_connection(334);
    `monitor_scoreboard_upstream_connection(335);
    `monitor_scoreboard_upstream_connection(336);
    `monitor_scoreboard_upstream_connection(337);
    `monitor_scoreboard_upstream_connection(338);
    `monitor_scoreboard_upstream_connection(339);
    `monitor_scoreboard_upstream_connection(340);
    `monitor_scoreboard_upstream_connection(341);
    `monitor_scoreboard_upstream_connection(342);
    `monitor_scoreboard_upstream_connection(343);
    `monitor_scoreboard_upstream_connection(344);
    `monitor_scoreboard_upstream_connection(345);
    `monitor_scoreboard_upstream_connection(346);
    `monitor_scoreboard_upstream_connection(347);
    `monitor_scoreboard_upstream_connection(348);
    `monitor_scoreboard_upstream_connection(349);
    `monitor_scoreboard_upstream_connection(350);
    `monitor_scoreboard_upstream_connection(351);
    `monitor_scoreboard_upstream_connection(352);
    `monitor_scoreboard_upstream_connection(353);
    `monitor_scoreboard_upstream_connection(354);
    `monitor_scoreboard_upstream_connection(355);
    `monitor_scoreboard_upstream_connection(356);
    `monitor_scoreboard_upstream_connection(357);
    `monitor_scoreboard_upstream_connection(358);
    `monitor_scoreboard_upstream_connection(359);
    `monitor_scoreboard_upstream_connection(360);
    `monitor_scoreboard_upstream_connection(361);
    `monitor_scoreboard_upstream_connection(362);
    `monitor_scoreboard_upstream_connection(363);
    `monitor_scoreboard_upstream_connection(364);
    `monitor_scoreboard_upstream_connection(365);
    `monitor_scoreboard_upstream_connection(366);
    `monitor_scoreboard_upstream_connection(367);
    `monitor_scoreboard_upstream_connection(368);
    `monitor_scoreboard_upstream_connection(369);
    `monitor_scoreboard_upstream_connection(370);
    `monitor_scoreboard_upstream_connection(371);
    `monitor_scoreboard_upstream_connection(372);
    `monitor_scoreboard_upstream_connection(373);
    `monitor_scoreboard_upstream_connection(374);
    `monitor_scoreboard_upstream_connection(375);
    `monitor_scoreboard_upstream_connection(376);
    `monitor_scoreboard_upstream_connection(377);
    `monitor_scoreboard_upstream_connection(378);
    `monitor_scoreboard_upstream_connection(379);
    `monitor_scoreboard_upstream_connection(380);
    `monitor_scoreboard_upstream_connection(381);
    `monitor_scoreboard_upstream_connection(382);
    `monitor_scoreboard_upstream_connection(383);
    `monitor_scoreboard_upstream_connection(384);
    `monitor_scoreboard_upstream_connection(385);
    `monitor_scoreboard_upstream_connection(386);
    `monitor_scoreboard_upstream_connection(387);
    `monitor_scoreboard_upstream_connection(388);
    `monitor_scoreboard_upstream_connection(389);
    `monitor_scoreboard_upstream_connection(390);
    `monitor_scoreboard_upstream_connection(391);
    `monitor_scoreboard_upstream_connection(392);
    `monitor_scoreboard_upstream_connection(393);
    `monitor_scoreboard_upstream_connection(394);
    `monitor_scoreboard_upstream_connection(395);
    `monitor_scoreboard_upstream_connection(396);
    `monitor_scoreboard_upstream_connection(397);
    `monitor_scoreboard_upstream_connection(398);
    `monitor_scoreboard_upstream_connection(399);
    `monitor_scoreboard_upstream_connection(400);
    `monitor_scoreboard_upstream_connection(401);
    `monitor_scoreboard_upstream_connection(402);
    `monitor_scoreboard_upstream_connection(403);
    `monitor_scoreboard_upstream_connection(404);
    `monitor_scoreboard_upstream_connection(405);
    `monitor_scoreboard_upstream_connection(406);
    `monitor_scoreboard_upstream_connection(407);
    `monitor_scoreboard_upstream_connection(408);
    `monitor_scoreboard_upstream_connection(409);
    `monitor_scoreboard_upstream_connection(410);
    `monitor_scoreboard_upstream_connection(411);
    `monitor_scoreboard_upstream_connection(412);
    `monitor_scoreboard_upstream_connection(413);
    `monitor_scoreboard_upstream_connection(414);
    `monitor_scoreboard_upstream_connection(415);
    `monitor_scoreboard_upstream_connection(416);
    `monitor_scoreboard_upstream_connection(417);
    `monitor_scoreboard_upstream_connection(418);
    `monitor_scoreboard_upstream_connection(419);
    `monitor_scoreboard_upstream_connection(420);
    `monitor_scoreboard_upstream_connection(421);
    `monitor_scoreboard_upstream_connection(422);
    `monitor_scoreboard_upstream_connection(423);
    `monitor_scoreboard_upstream_connection(424);
    `monitor_scoreboard_upstream_connection(425);
    `monitor_scoreboard_upstream_connection(426);
    `monitor_scoreboard_upstream_connection(427);
    `monitor_scoreboard_upstream_connection(428);
    `monitor_scoreboard_upstream_connection(429);
    `monitor_scoreboard_upstream_connection(430);
    `monitor_scoreboard_upstream_connection(431);
    `monitor_scoreboard_upstream_connection(432);
    `monitor_scoreboard_upstream_connection(433);
    `monitor_scoreboard_upstream_connection(434);
    `monitor_scoreboard_upstream_connection(435);
    `monitor_scoreboard_upstream_connection(436);
    `monitor_scoreboard_upstream_connection(437);
    `monitor_scoreboard_upstream_connection(438);
    `monitor_scoreboard_upstream_connection(439);
    `monitor_scoreboard_upstream_connection(440);
    `monitor_scoreboard_upstream_connection(441);
    `monitor_scoreboard_upstream_connection(442);
    `monitor_scoreboard_upstream_connection(443);
    `monitor_scoreboard_upstream_connection(444);
    `monitor_scoreboard_upstream_connection(445);
    `monitor_scoreboard_upstream_connection(446);
    `monitor_scoreboard_upstream_connection(447);
    `monitor_scoreboard_upstream_connection(448);
    `monitor_scoreboard_upstream_connection(449);
    `monitor_scoreboard_upstream_connection_TB4(0,450,0);
    `monitor_scoreboard_upstream_connection_TB4(0,451,1);
    `monitor_scoreboard_upstream_connection_TB4(0,452,2);
    `monitor_scoreboard_upstream_connection_TB4(0,453,3);
    `monitor_scoreboard_upstream_connection_TB4(0,454,4);
    `monitor_scoreboard_upstream_connection_TB4(0,455,5);
    `monitor_scoreboard_upstream_connection_TB4(0,456,6);
    `monitor_scoreboard_upstream_connection_TB4(0,457,7);
    `monitor_scoreboard_upstream_connection_TB4(0,458,8);
    `monitor_scoreboard_upstream_connection_TB4(0,459,9);
    `monitor_scoreboard_upstream_connection_TB4(0,460,10);
    `monitor_scoreboard_upstream_connection_TB4(0,461,11);
    `monitor_scoreboard_upstream_connection_TB4(0,462,12);
    `monitor_scoreboard_upstream_connection_TB4(0,463,13);
    `monitor_scoreboard_upstream_connection_TB4(0,464,14);
    `monitor_scoreboard_upstream_connection_TB4(0,465,15);
    `monitor_scoreboard_upstream_connection_TB4(0,466,16);
    `monitor_scoreboard_upstream_connection_TB4(0,467,17);
    `monitor_scoreboard_upstream_connection_TB4(0,468,18);
    `monitor_scoreboard_upstream_connection_TB4(0,469,19);
    `monitor_scoreboard_upstream_connection_TB4(0,470,20);
    `monitor_scoreboard_upstream_connection_TB4(0,471,21);
    `monitor_scoreboard_upstream_connection_TB4(0,472,22);
    `monitor_scoreboard_upstream_connection_TB4(0,473,23);
    `monitor_scoreboard_upstream_connection_TB4(0,474,24);
    `monitor_scoreboard_upstream_connection_TB4(0,475,25);
    `monitor_scoreboard_upstream_connection_TB4(0,476,26);
    `monitor_scoreboard_upstream_connection_TB4(0,477,27);
    `monitor_scoreboard_upstream_connection_TB4(0,478,28);
    `monitor_scoreboard_upstream_connection_TB4(0,479,29);
    `monitor_scoreboard_upstream_connection_TB4(0,480,30);
    `monitor_scoreboard_upstream_connection_TB4(0,481,31);
    `monitor_scoreboard_upstream_connection_TB4(0,482,32);
    `monitor_scoreboard_upstream_connection_TB4(0,483,33);
    `monitor_scoreboard_upstream_connection_TB4(0,484,34);
    `monitor_scoreboard_upstream_connection_TB4(0,485,35);
    `monitor_scoreboard_upstream_connection_TB4(0,486,36);
    `monitor_scoreboard_upstream_connection_TB4(0,487,37);
    `monitor_scoreboard_upstream_connection_TB4(0,488,38);
    `monitor_scoreboard_upstream_connection_TB4(0,489,39);
    `monitor_scoreboard_upstream_connection_TB4(0,490,40);
    `monitor_scoreboard_upstream_connection_TB4(0,491,41);
    `monitor_scoreboard_upstream_connection_TB4(0,492,42);
    `monitor_scoreboard_upstream_connection_TB4(0,493,43);
    `monitor_scoreboard_upstream_connection_TB4(0,494,44);
    `monitor_scoreboard_upstream_connection_TB4(0,495,45);
    `monitor_scoreboard_upstream_connection_TB4(0,496,46);
    `monitor_scoreboard_upstream_connection_TB4(0,497,47);
    `monitor_scoreboard_upstream_connection_TB4(0,498,48);
    `monitor_scoreboard_upstream_connection_TB4(0,499,49);
    `monitor_scoreboard_upstream_connection_TB4(0,500,50);
    `monitor_scoreboard_upstream_connection_TB4(0,501,51);
    `monitor_scoreboard_upstream_connection_TB4(0,502,52);
    `monitor_scoreboard_upstream_connection_TB4(0,503,53);
    `monitor_scoreboard_upstream_connection_TB4(0,504,54);
    `monitor_scoreboard_upstream_connection_TB4(0,505,55);
    `monitor_scoreboard_upstream_connection_TB4(0,506,56);
    `monitor_scoreboard_upstream_connection_TB4(0,507,57);
    `monitor_scoreboard_upstream_connection_TB4(0,508,58);
    `monitor_scoreboard_upstream_connection_TB4(0,509,59);
    `monitor_scoreboard_upstream_connection_TB4(0,510,60);
    `monitor_scoreboard_upstream_connection_TB4(0,511,61);
    `monitor_scoreboard_upstream_connection_TB4(0,512,62);
    `monitor_scoreboard_upstream_connection_TB4(0,513,63);
    `monitor_scoreboard_upstream_connection_TB4(0,514,64);
    `monitor_scoreboard_upstream_connection_TB4(0,515,65);
    `monitor_scoreboard_upstream_connection_TB4(0,516,66);
    `monitor_scoreboard_upstream_connection_TB4(0,517,67);
    `monitor_scoreboard_upstream_connection_TB4(0,518,68);
    `monitor_scoreboard_upstream_connection_TB4(0,519,69);
    `monitor_scoreboard_upstream_connection_TB4(0,520,70);
    `monitor_scoreboard_upstream_connection_TB4(0,521,71);
    `monitor_scoreboard_upstream_connection_TB4(0,522,72);
    `monitor_scoreboard_upstream_connection_TB4(0,523,73);
    `monitor_scoreboard_upstream_connection_TB4(0,524,74);
    `monitor_scoreboard_upstream_connection_TB4(0,525,75);
    `monitor_scoreboard_upstream_connection_TB4(0,526,76);
    `monitor_scoreboard_upstream_connection_TB4(0,527,77);
    `monitor_scoreboard_upstream_connection_TB4(0,528,78);
    `monitor_scoreboard_upstream_connection_TB4(0,529,79);
    `monitor_scoreboard_upstream_connection_TB4(0,530,80);
    `monitor_scoreboard_upstream_connection_TB4(0,531,81);
    `monitor_scoreboard_upstream_connection_TB4(0,532,82);
    `monitor_scoreboard_upstream_connection_TB4(0,533,83);
    `monitor_scoreboard_upstream_connection_TB4(0,534,84);
    `monitor_scoreboard_upstream_connection_TB4(0,535,85);
    `monitor_scoreboard_upstream_connection_TB4(0,536,86);
    `monitor_scoreboard_upstream_connection_TB4(0,537,87);
    `monitor_scoreboard_upstream_connection_TB4(0,538,88);
    `monitor_scoreboard_upstream_connection_TB4(0,539,89);
    `monitor_scoreboard_upstream_connection_TB4(0,540,90);
    `monitor_scoreboard_upstream_connection_TB4(0,541,91);
    `monitor_scoreboard_upstream_connection_TB4(0,542,92);
    `monitor_scoreboard_upstream_connection_TB4(0,543,93);
    `monitor_scoreboard_upstream_connection_TB4(0,544,94);
    `monitor_scoreboard_upstream_connection_TB4(0,545,95);
    `monitor_scoreboard_upstream_connection_TB4(0,546,96);
    `monitor_scoreboard_upstream_connection_TB4(0,547,97);
    `monitor_scoreboard_upstream_connection_TB4(0,548,98);
    `monitor_scoreboard_upstream_connection_TB4(0,549,99);
    `monitor_scoreboard_upstream_connection_TB4(0,550,100);
    `monitor_scoreboard_upstream_connection_TB4(0,551,101);
    `monitor_scoreboard_upstream_connection_TB4(0,552,102);
    `monitor_scoreboard_upstream_connection_TB4(0,553,103);
    `monitor_scoreboard_upstream_connection_TB4(0,554,104);
    `monitor_scoreboard_upstream_connection_TB4(0,555,105);
    `monitor_scoreboard_upstream_connection_TB4(0,556,106);
    `monitor_scoreboard_upstream_connection_TB4(0,557,107);
    `monitor_scoreboard_upstream_connection_TB4(0,558,108);
    `monitor_scoreboard_upstream_connection_TB4(0,559,109);
    `monitor_scoreboard_upstream_connection_TB4(0,560,110);
    `monitor_scoreboard_upstream_connection_TB4(0,561,111);
    `monitor_scoreboard_upstream_connection_TB4(0,562,112);
    `monitor_scoreboard_upstream_connection_TB4(0,563,113);
    `monitor_scoreboard_upstream_connection_TB4(0,564,114);
    `monitor_scoreboard_upstream_connection_TB4(0,565,115);
    `monitor_scoreboard_upstream_connection_TB4(0,566,116);
    `monitor_scoreboard_upstream_connection_TB4(0,567,117);
    `monitor_scoreboard_upstream_connection_TB4(0,568,118);
    `monitor_scoreboard_upstream_connection_TB4(0,569,119);
    `monitor_scoreboard_upstream_connection_TB4(0,570,120);
    `monitor_scoreboard_upstream_connection_TB4(0,571,121);
    `monitor_scoreboard_upstream_connection_TB4(0,572,122);
    `monitor_scoreboard_upstream_connection_TB4(0,573,123);
    `monitor_scoreboard_upstream_connection_TB4(0,574,124);
    `monitor_scoreboard_upstream_connection_TB4(0,575,125);
    `monitor_scoreboard_upstream_connection_TB4(0,576,126);
    `monitor_scoreboard_upstream_connection_TB4(0,577,127);
    `monitor_scoreboard_upstream_connection_TB4(0,578,128);
    `monitor_scoreboard_upstream_connection_TB4(0,579,129);
    `monitor_scoreboard_upstream_connection_TB4(0,580,130);
    `monitor_scoreboard_upstream_connection_TB4(0,581,131);
    `monitor_scoreboard_upstream_connection_TB4(0,582,132);
    `monitor_scoreboard_upstream_connection_TB4(0,583,133);
    `monitor_scoreboard_upstream_connection_TB4(0,584,134);
    `monitor_scoreboard_upstream_connection_TB4(0,585,135);
    `monitor_scoreboard_upstream_connection_TB4(0,586,136);
    `monitor_scoreboard_upstream_connection_TB4(0,587,137);
    `monitor_scoreboard_upstream_connection_TB4(0,588,138);
    `monitor_scoreboard_upstream_connection_TB4(0,589,139);
    `monitor_scoreboard_upstream_connection_TB4(0,590,140);
    `monitor_scoreboard_upstream_connection_TB4(0,591,141);
    `monitor_scoreboard_upstream_connection_TB4(0,592,142);
    `monitor_scoreboard_upstream_connection_TB4(0,593,143);
    `monitor_scoreboard_upstream_connection_TB4(0,594,144);
    `monitor_scoreboard_upstream_connection_TB4(0,595,145);
    `monitor_scoreboard_upstream_connection_TB4(0,596,146);
    `monitor_scoreboard_upstream_connection_TB4(0,597,147);
    `monitor_scoreboard_upstream_connection_TB4(0,598,148);
    `monitor_scoreboard_upstream_connection_TB4(0,599,149);
    `monitor_scoreboard_upstream_connection_TB4(0,600,150);
    `monitor_scoreboard_upstream_connection_TB4(0,601,151);
    `monitor_scoreboard_upstream_connection_TB4(0,602,152);
    `monitor_scoreboard_upstream_connection_TB4(0,603,153);
    `monitor_scoreboard_upstream_connection_TB4(0,604,154);
    `monitor_scoreboard_upstream_connection_TB4(0,605,155);
    `monitor_scoreboard_upstream_connection_TB4(0,606,156);
    `monitor_scoreboard_upstream_connection_TB4(0,607,157);
    `monitor_scoreboard_upstream_connection_TB4(0,608,158);
    `monitor_scoreboard_upstream_connection_TB4(0,609,159);
    `monitor_scoreboard_upstream_connection_TB4(0,610,160);
    `monitor_scoreboard_upstream_connection_TB4(0,611,161);
    `monitor_scoreboard_upstream_connection_TB4(0,612,162);
    `monitor_scoreboard_upstream_connection_TB4(0,613,163);
    `monitor_scoreboard_upstream_connection_TB4(0,614,164);
    `monitor_scoreboard_upstream_connection_TB4(0,615,165);
    `monitor_scoreboard_upstream_connection_TB4(0,616,166);
    `monitor_scoreboard_upstream_connection_TB4(0,617,167);
    `monitor_scoreboard_upstream_connection_TB4(0,618,168);
    `monitor_scoreboard_upstream_connection_TB4(0,619,169);
    `monitor_scoreboard_upstream_connection_TB4(0,620,170);
    `monitor_scoreboard_upstream_connection_TB4(0,621,171);
    `monitor_scoreboard_upstream_connection_TB4(0,622,172);
    `monitor_scoreboard_upstream_connection_TB4(0,623,173);
    `monitor_scoreboard_upstream_connection_TB4(0,624,174);
    `monitor_scoreboard_upstream_connection_TB4(0,625,175);
    `monitor_scoreboard_upstream_connection_TB4(0,626,176);
    `monitor_scoreboard_upstream_connection_TB4(0,627,177);
    `monitor_scoreboard_upstream_connection_TB4(0,628,178);
    `monitor_scoreboard_upstream_connection_TB4(0,629,179);
    `monitor_scoreboard_upstream_connection_TB4(0,630,180);
    `monitor_scoreboard_upstream_connection_TB4(0,631,181);
    `monitor_scoreboard_upstream_connection_TB4(0,632,182);
    `monitor_scoreboard_upstream_connection_TB4(0,633,183);
    `monitor_scoreboard_upstream_connection_TB4(0,634,184);
    `monitor_scoreboard_upstream_connection_TB4(0,635,185);
    `monitor_scoreboard_upstream_connection_TB4(0,636,186);
    `monitor_scoreboard_upstream_connection_TB4(0,637,187);
    `monitor_scoreboard_upstream_connection_TB4(0,638,188);
    `monitor_scoreboard_upstream_connection_TB4(0,639,189);
    `monitor_scoreboard_upstream_connection_TB4(0,640,190);
    `monitor_scoreboard_upstream_connection_TB4(0,641,191);
    `monitor_scoreboard_upstream_connection_TB4(0,642,192);
    `monitor_scoreboard_upstream_connection_TB4(0,643,193);
    `monitor_scoreboard_upstream_connection_TB4(0,644,194);
    `monitor_scoreboard_upstream_connection_TB4(0,645,195);
    `monitor_scoreboard_upstream_connection_TB4(0,646,196);
    `monitor_scoreboard_upstream_connection_TB4(0,647,197);
    `monitor_scoreboard_upstream_connection_TB4(0,648,198);
    `monitor_scoreboard_upstream_connection_TB4(0,649,199);
    `monitor_scoreboard_upstream_connection_TB4(0,650,200);
    `monitor_scoreboard_upstream_connection_TB4(0,651,201);
    `monitor_scoreboard_upstream_connection_TB4(0,652,202);
    `monitor_scoreboard_upstream_connection_TB4(0,653,203);
    `monitor_scoreboard_upstream_connection_TB4(0,654,204);
    `monitor_scoreboard_upstream_connection_TB4(0,655,205);
    `monitor_scoreboard_upstream_connection_TB4(0,656,206);
    `monitor_scoreboard_upstream_connection_TB4(0,657,207);
    `monitor_scoreboard_upstream_connection_TB4(0,658,208);
    `monitor_scoreboard_upstream_connection_TB4(0,659,209);
    `monitor_scoreboard_upstream_connection_TB4(0,660,210);
    `monitor_scoreboard_upstream_connection_TB4(0,661,211);
    `monitor_scoreboard_upstream_connection_TB4(0,662,212);
    `monitor_scoreboard_upstream_connection_TB4(0,663,213);
    `monitor_scoreboard_upstream_connection_TB4(0,664,214);
    `monitor_scoreboard_upstream_connection_TB4(0,665,215);
    `monitor_scoreboard_upstream_connection_TB4(0,666,216);
    `monitor_scoreboard_upstream_connection_TB4(0,667,217);
    `monitor_scoreboard_upstream_connection_TB4(0,668,218);
    `monitor_scoreboard_upstream_connection_TB4(0,669,219);
    `monitor_scoreboard_upstream_connection_TB4(0,670,220);
    `monitor_scoreboard_upstream_connection_TB4(0,671,221);
    `monitor_scoreboard_upstream_connection_TB4(0,672,222);
    `monitor_scoreboard_upstream_connection_TB4(0,673,223);
    `monitor_scoreboard_upstream_connection_TB4(0,674,224);
    `monitor_scoreboard_upstream_connection_TB4(0,675,225);
    `monitor_scoreboard_upstream_connection_TB4(0,676,226);
    `monitor_scoreboard_upstream_connection_TB4(0,677,227);
    `monitor_scoreboard_upstream_connection_TB4(0,678,228);
    `monitor_scoreboard_upstream_connection_TB4(0,679,229);
    `monitor_scoreboard_upstream_connection_TB4(0,680,230);
    `monitor_scoreboard_upstream_connection_TB4(0,681,231);
    `monitor_scoreboard_upstream_connection_TB4(0,682,232);
    `monitor_scoreboard_upstream_connection_TB4(0,683,233);
    `monitor_scoreboard_upstream_connection_TB4(0,684,234);
    `monitor_scoreboard_upstream_connection_TB4(0,685,235);
    `monitor_scoreboard_upstream_connection_TB4(0,686,236);
    `monitor_scoreboard_upstream_connection_TB4(0,687,237);
    `monitor_scoreboard_upstream_connection_TB4(0,688,238);
    `monitor_scoreboard_upstream_connection_TB4(0,689,239);
    `monitor_scoreboard_upstream_connection_TB4(0,690,240);
    `monitor_scoreboard_upstream_connection_TB4(0,691,241);
    `monitor_scoreboard_upstream_connection_TB4(0,692,242);
    `monitor_scoreboard_upstream_connection_TB4(0,693,243);
    `monitor_scoreboard_upstream_connection_TB4(0,694,244);
    `monitor_scoreboard_upstream_connection_TB4(0,695,245);
    `monitor_scoreboard_upstream_connection_TB4(0,696,246);
    `monitor_scoreboard_upstream_connection_TB4(0,697,247);
    `monitor_scoreboard_upstream_connection_TB4(0,698,248);
    `monitor_scoreboard_upstream_connection_TB4(0,699,249);
    `monitor_scoreboard_upstream_connection_TB4(0,700,250);
    `monitor_scoreboard_upstream_connection_TB4(0,701,251);
    `monitor_scoreboard_upstream_connection_TB4(0,702,252);
    `monitor_scoreboard_upstream_connection_TB4(0,703,253);
    `monitor_scoreboard_upstream_connection_TB4(0,704,254);
    `monitor_scoreboard_upstream_connection_TB4(0,705,255);
    `monitor_scoreboard_upstream_connection_TB4(0,706,256);
    `monitor_scoreboard_upstream_connection_TB4(0,707,257);
    `monitor_scoreboard_upstream_connection_TB4(0,708,258);
    `monitor_scoreboard_upstream_connection_TB4(0,709,259);
    `monitor_scoreboard_upstream_connection_TB4(0,710,260);
    `monitor_scoreboard_upstream_connection_TB4(0,711,261);
    `monitor_scoreboard_upstream_connection_TB4(0,712,262);
    `monitor_scoreboard_upstream_connection_TB4(0,713,263);
    `monitor_scoreboard_upstream_connection_TB4(0,714,264);
    `monitor_scoreboard_upstream_connection_TB4(0,715,265);
    `monitor_scoreboard_upstream_connection_TB4(0,716,266);
    `monitor_scoreboard_upstream_connection_TB4(0,717,267);
    `monitor_scoreboard_upstream_connection_TB4(0,718,268);
    `monitor_scoreboard_upstream_connection_TB4(0,719,269);
    `monitor_scoreboard_upstream_connection_TB4(0,720,270);
    `monitor_scoreboard_upstream_connection_TB4(0,721,271);
    `monitor_scoreboard_upstream_connection_TB4(0,722,272);
    `monitor_scoreboard_upstream_connection_TB4(0,723,273);
    `monitor_scoreboard_upstream_connection_TB4(0,724,274);
    `monitor_scoreboard_upstream_connection_TB4(0,725,275);
    `monitor_scoreboard_upstream_connection_TB4(0,726,276);
    `monitor_scoreboard_upstream_connection_TB4(0,727,277);
    `monitor_scoreboard_upstream_connection_TB4(0,728,278);
    `monitor_scoreboard_upstream_connection_TB4(0,729,279);
    `monitor_scoreboard_upstream_connection_TB4(0,730,280);
    `monitor_scoreboard_upstream_connection_TB4(0,731,281);
    `monitor_scoreboard_upstream_connection_TB4(0,732,282);
    `monitor_scoreboard_upstream_connection_TB4(0,733,283);
    `monitor_scoreboard_upstream_connection_TB4(0,734,284);
    `monitor_scoreboard_upstream_connection_TB4(0,735,285);
    `monitor_scoreboard_upstream_connection_TB4(0,736,286);
    `monitor_scoreboard_upstream_connection_TB4(0,737,287);
    `monitor_scoreboard_upstream_connection_TB4(0,738,288);
    `monitor_scoreboard_upstream_connection_TB4(0,739,289);
    `monitor_scoreboard_upstream_connection_TB4(0,740,290);
    `monitor_scoreboard_upstream_connection_TB4(0,741,291);
    `monitor_scoreboard_upstream_connection_TB4(0,742,292);
    `monitor_scoreboard_upstream_connection_TB4(0,743,293);
    `monitor_scoreboard_upstream_connection_TB4(0,744,294);
    `monitor_scoreboard_upstream_connection_TB4(0,745,295);
    `monitor_scoreboard_upstream_connection_TB4(0,746,296);
    `monitor_scoreboard_upstream_connection_TB4(0,747,297);
    `monitor_scoreboard_upstream_connection_TB4(0,748,298);
    `monitor_scoreboard_upstream_connection_TB4(0,749,299);
    `monitor_scoreboard_upstream_connection_TB4(0,750,300);
    `monitor_scoreboard_upstream_connection_TB4(0,751,301);
    `monitor_scoreboard_upstream_connection_TB4(0,752,302);
    `monitor_scoreboard_upstream_connection_TB4(0,753,303);
    `monitor_scoreboard_upstream_connection_TB4(0,754,304);
    `monitor_scoreboard_upstream_connection_TB4(0,755,305);
    `monitor_scoreboard_upstream_connection_TB4(0,756,306);
    `monitor_scoreboard_upstream_connection_TB4(0,757,307);
    `monitor_scoreboard_upstream_connection_TB4(0,758,308);
    `monitor_scoreboard_upstream_connection_TB4(0,759,309);
    `monitor_scoreboard_upstream_connection_TB4(0,760,310);
    `monitor_scoreboard_upstream_connection_TB4(0,761,311);
    `monitor_scoreboard_upstream_connection_TB4(0,762,312);
    `monitor_scoreboard_upstream_connection_TB4(0,763,313);
    `monitor_scoreboard_upstream_connection_TB4(0,764,314);
    `monitor_scoreboard_upstream_connection_TB4(0,765,315);
    `monitor_scoreboard_upstream_connection_TB4(0,766,316);
    `monitor_scoreboard_upstream_connection_TB4(0,767,317);
    `monitor_scoreboard_upstream_connection_TB4(0,768,318);
    `monitor_scoreboard_upstream_connection_TB4(0,769,319);
    `monitor_scoreboard_upstream_connection_TB4(0,770,320);
    `monitor_scoreboard_upstream_connection_TB4(0,771,321);
    `monitor_scoreboard_upstream_connection_TB4(0,772,322);
    `monitor_scoreboard_upstream_connection_TB4(0,773,323);
    `monitor_scoreboard_upstream_connection_TB4(0,774,324);
    `monitor_scoreboard_upstream_connection_TB4(0,775,325);
    `monitor_scoreboard_upstream_connection_TB4(0,776,326);
    `monitor_scoreboard_upstream_connection_TB4(0,777,327);
    `monitor_scoreboard_upstream_connection_TB4(0,778,328);
    `monitor_scoreboard_upstream_connection_TB4(0,779,329);
    `monitor_scoreboard_upstream_connection_TB4(0,780,330);
    `monitor_scoreboard_upstream_connection_TB4(0,781,331);
    `monitor_scoreboard_upstream_connection_TB4(0,782,332);
    `monitor_scoreboard_upstream_connection_TB4(0,783,333);
    `monitor_scoreboard_upstream_connection_TB4(0,784,334);
    `monitor_scoreboard_upstream_connection_TB4(0,785,335);
    `monitor_scoreboard_upstream_connection_TB4(0,786,336);
    `monitor_scoreboard_upstream_connection_TB4(0,787,337);
    `monitor_scoreboard_upstream_connection_TB4(0,788,338);
    `monitor_scoreboard_upstream_connection_TB4(0,789,339);
    `monitor_scoreboard_upstream_connection_TB4(0,790,340);
    `monitor_scoreboard_upstream_connection_TB4(0,791,341);
    `monitor_scoreboard_upstream_connection_TB4(0,792,342);
    `monitor_scoreboard_upstream_connection_TB4(0,793,343);
    `monitor_scoreboard_upstream_connection_TB4(0,794,344);
    `monitor_scoreboard_upstream_connection_TB4(0,795,345);
    `monitor_scoreboard_upstream_connection_TB4(0,796,346);
    `monitor_scoreboard_upstream_connection_TB4(0,797,347);
    `monitor_scoreboard_upstream_connection_TB4(0,798,348);
    `monitor_scoreboard_upstream_connection_TB4(0,799,349);
    `monitor_scoreboard_upstream_connection_TB4(0,800,350);
    `monitor_scoreboard_upstream_connection_TB4(0,801,351);
    `monitor_scoreboard_upstream_connection_TB4(0,802,352);
    `monitor_scoreboard_upstream_connection_TB4(0,803,353);
    `monitor_scoreboard_upstream_connection_TB4(0,804,354);
    `monitor_scoreboard_upstream_connection_TB4(0,805,355);
    `monitor_scoreboard_upstream_connection_TB4(0,806,356);
    `monitor_scoreboard_upstream_connection_TB4(0,807,357);
    `monitor_scoreboard_upstream_connection_TB4(0,808,358);
    `monitor_scoreboard_upstream_connection_TB4(0,809,359);
    `monitor_scoreboard_upstream_connection_TB4(0,810,360);
    `monitor_scoreboard_upstream_connection_TB4(0,811,361);
    `monitor_scoreboard_upstream_connection_TB4(0,812,362);
    `monitor_scoreboard_upstream_connection_TB4(0,813,363);
    `monitor_scoreboard_upstream_connection_TB4(0,814,364);
    `monitor_scoreboard_upstream_connection_TB4(0,815,365);
    `monitor_scoreboard_upstream_connection_TB4(0,816,366);
    `monitor_scoreboard_upstream_connection_TB4(0,817,367);
    `monitor_scoreboard_upstream_connection_TB4(0,818,368);
    `monitor_scoreboard_upstream_connection_TB4(0,819,369);
    `monitor_scoreboard_upstream_connection_TB4(0,820,370);
    `monitor_scoreboard_upstream_connection_TB4(0,821,371);
    `monitor_scoreboard_upstream_connection_TB4(0,822,372);
    `monitor_scoreboard_upstream_connection_TB4(0,823,373);
    `monitor_scoreboard_upstream_connection_TB4(0,824,374);
    `monitor_scoreboard_upstream_connection_TB4(0,825,375);
    `monitor_scoreboard_upstream_connection_TB4(0,826,376);
    `monitor_scoreboard_upstream_connection_TB4(0,827,377);
    `monitor_scoreboard_upstream_connection_TB4(0,828,378);
    `monitor_scoreboard_upstream_connection_TB4(0,829,379);
    `monitor_scoreboard_upstream_connection_TB4(0,830,380);
    `monitor_scoreboard_upstream_connection_TB4(0,831,381);
    `monitor_scoreboard_upstream_connection_TB4(0,832,382);
    `monitor_scoreboard_upstream_connection_TB4(0,833,383);
    `monitor_scoreboard_upstream_connection_TB4(0,834,384);
    `monitor_scoreboard_upstream_connection_TB4(0,835,385);
    `monitor_scoreboard_upstream_connection_TB4(0,836,386);
    `monitor_scoreboard_upstream_connection_TB4(0,837,387);
    `monitor_scoreboard_upstream_connection_TB4(0,838,388);
    `monitor_scoreboard_upstream_connection_TB4(0,839,389);
    `monitor_scoreboard_upstream_connection_TB4(0,840,390);
    `monitor_scoreboard_upstream_connection_TB4(0,841,391);
    `monitor_scoreboard_upstream_connection_TB4(0,842,392);
    `monitor_scoreboard_upstream_connection_TB4(0,843,393);
    `monitor_scoreboard_upstream_connection_TB4(0,844,394);
    `monitor_scoreboard_upstream_connection_TB4(0,845,395);
    `monitor_scoreboard_upstream_connection_TB4(0,846,396);
    `monitor_scoreboard_upstream_connection_TB4(0,847,397);
    `monitor_scoreboard_upstream_connection_TB4(0,848,398);
    `monitor_scoreboard_upstream_connection_TB4(0,849,399);
    `monitor_scoreboard_upstream_connection_TB4(0,850,400);
    `monitor_scoreboard_upstream_connection_TB4(0,851,401);
    `monitor_scoreboard_upstream_connection_TB4(0,852,402);
    `monitor_scoreboard_upstream_connection_TB4(0,853,403);
    `monitor_scoreboard_upstream_connection_TB4(0,854,404);
    `monitor_scoreboard_upstream_connection_TB4(0,855,405);
    `monitor_scoreboard_upstream_connection_TB4(0,856,406);
    `monitor_scoreboard_upstream_connection_TB4(0,857,407);
    `monitor_scoreboard_upstream_connection_TB4(0,858,408);
    `monitor_scoreboard_upstream_connection_TB4(0,859,409);
    `monitor_scoreboard_upstream_connection_TB4(0,860,410);
    `monitor_scoreboard_upstream_connection_TB4(0,861,411);
    `monitor_scoreboard_upstream_connection_TB4(0,862,412);
    `monitor_scoreboard_upstream_connection_TB4(0,863,413);
    `monitor_scoreboard_upstream_connection_TB4(0,864,414);
    `monitor_scoreboard_upstream_connection_TB4(0,865,415);
    `monitor_scoreboard_upstream_connection_TB4(0,866,416);
    `monitor_scoreboard_upstream_connection_TB4(0,867,417);
    `monitor_scoreboard_upstream_connection_TB4(0,868,418);
    `monitor_scoreboard_upstream_connection_TB4(0,869,419);
    `monitor_scoreboard_upstream_connection_TB4(0,870,420);
    `monitor_scoreboard_upstream_connection_TB4(0,871,421);
    `monitor_scoreboard_upstream_connection_TB4(0,872,422);
    `monitor_scoreboard_upstream_connection_TB4(0,873,423);
    `monitor_scoreboard_upstream_connection_TB4(0,874,424);
    `monitor_scoreboard_upstream_connection_TB4(0,875,425);
    `monitor_scoreboard_upstream_connection_TB4(0,876,426);
    `monitor_scoreboard_upstream_connection_TB4(0,877,427);
    `monitor_scoreboard_upstream_connection_TB4(0,878,428);
    `monitor_scoreboard_upstream_connection_TB4(0,879,429);
    `monitor_scoreboard_upstream_connection_TB4(0,880,430);
    `monitor_scoreboard_upstream_connection_TB4(0,881,431);
    `monitor_scoreboard_upstream_connection_TB4(0,882,432);
    `monitor_scoreboard_upstream_connection_TB4(0,883,433);
    `monitor_scoreboard_upstream_connection_TB4(0,884,434);
    `monitor_scoreboard_upstream_connection_TB4(0,885,435);
    `monitor_scoreboard_upstream_connection_TB4(0,886,436);
    `monitor_scoreboard_upstream_connection_TB4(0,887,437);
    `monitor_scoreboard_upstream_connection_TB4(0,888,438);
    `monitor_scoreboard_upstream_connection_TB4(0,889,439);
    `monitor_scoreboard_upstream_connection_TB4(0,890,440);
    `monitor_scoreboard_upstream_connection_TB4(0,891,441);
    `monitor_scoreboard_upstream_connection_TB4(0,892,442);
    `monitor_scoreboard_upstream_connection_TB4(0,893,443);
    `monitor_scoreboard_upstream_connection_TB4(0,894,444);
    `monitor_scoreboard_upstream_connection_TB4(0,895,445);
    `monitor_scoreboard_upstream_connection_TB4(0,896,446);
    `monitor_scoreboard_upstream_connection_TB4(0,897,447);
    `monitor_scoreboard_upstream_connection_TB4(0,898,448);
    `monitor_scoreboard_upstream_connection_TB4(0,899,449);
    `monitor_scoreboard_upstream_connection_TB4(1,900,0);
    `monitor_scoreboard_upstream_connection_TB4(1,901,1);
    `monitor_scoreboard_upstream_connection_TB4(1,902,2);
    `monitor_scoreboard_upstream_connection_TB4(1,903,3);
    `monitor_scoreboard_upstream_connection_TB4(1,904,4);
    `monitor_scoreboard_upstream_connection_TB4(1,905,5);
    `monitor_scoreboard_upstream_connection_TB4(1,906,6);
    `monitor_scoreboard_upstream_connection_TB4(1,907,7);
    `monitor_scoreboard_upstream_connection_TB4(1,908,8);
    `monitor_scoreboard_upstream_connection_TB4(1,909,9);
    `monitor_scoreboard_upstream_connection_TB4(1,910,10);
    `monitor_scoreboard_upstream_connection_TB4(1,911,11);
    `monitor_scoreboard_upstream_connection_TB4(1,912,12);
    `monitor_scoreboard_upstream_connection_TB4(1,913,13);
    `monitor_scoreboard_upstream_connection_TB4(1,914,14);
    `monitor_scoreboard_upstream_connection_TB4(1,915,15);
    `monitor_scoreboard_upstream_connection_TB4(1,916,16);
    `monitor_scoreboard_upstream_connection_TB4(1,917,17);
    `monitor_scoreboard_upstream_connection_TB4(1,918,18);
    `monitor_scoreboard_upstream_connection_TB4(1,919,19);
    `monitor_scoreboard_upstream_connection_TB4(1,920,20);
    `monitor_scoreboard_upstream_connection_TB4(1,921,21);
    `monitor_scoreboard_upstream_connection_TB4(1,922,22);
    `monitor_scoreboard_upstream_connection_TB4(1,923,23);
    `monitor_scoreboard_upstream_connection_TB4(1,924,24);
    `monitor_scoreboard_upstream_connection_TB4(1,925,25);
    `monitor_scoreboard_upstream_connection_TB4(1,926,26);
    `monitor_scoreboard_upstream_connection_TB4(1,927,27);
    `monitor_scoreboard_upstream_connection_TB4(1,928,28);
    `monitor_scoreboard_upstream_connection_TB4(1,929,29);
    `monitor_scoreboard_upstream_connection_TB4(1,930,30);
    `monitor_scoreboard_upstream_connection_TB4(1,931,31);
    `monitor_scoreboard_upstream_connection_TB4(1,932,32);
    `monitor_scoreboard_upstream_connection_TB4(1,933,33);
    `monitor_scoreboard_upstream_connection_TB4(1,934,34);
    `monitor_scoreboard_upstream_connection_TB4(1,935,35);
    `monitor_scoreboard_upstream_connection_TB4(1,936,36);
    `monitor_scoreboard_upstream_connection_TB4(1,937,37);
    `monitor_scoreboard_upstream_connection_TB4(1,938,38);
    `monitor_scoreboard_upstream_connection_TB4(1,939,39);
    `monitor_scoreboard_upstream_connection_TB4(1,940,40);
    `monitor_scoreboard_upstream_connection_TB4(1,941,41);
    `monitor_scoreboard_upstream_connection_TB4(1,942,42);
    `monitor_scoreboard_upstream_connection_TB4(1,943,43);
    `monitor_scoreboard_upstream_connection_TB4(1,944,44);
    `monitor_scoreboard_upstream_connection_TB4(1,945,45);
    `monitor_scoreboard_upstream_connection_TB4(1,946,46);
    `monitor_scoreboard_upstream_connection_TB4(1,947,47);
    `monitor_scoreboard_upstream_connection_TB4(1,948,48);
    `monitor_scoreboard_upstream_connection_TB4(1,949,49);
    `monitor_scoreboard_upstream_connection_TB4(1,950,50);
    `monitor_scoreboard_upstream_connection_TB4(1,951,51);
    `monitor_scoreboard_upstream_connection_TB4(1,952,52);
    `monitor_scoreboard_upstream_connection_TB4(1,953,53);
    `monitor_scoreboard_upstream_connection_TB4(1,954,54);
    `monitor_scoreboard_upstream_connection_TB4(1,955,55);
    `monitor_scoreboard_upstream_connection_TB4(1,956,56);
    `monitor_scoreboard_upstream_connection_TB4(1,957,57);
    `monitor_scoreboard_upstream_connection_TB4(1,958,58);
    `monitor_scoreboard_upstream_connection_TB4(1,959,59);
    `monitor_scoreboard_upstream_connection_TB4(1,960,60);
    `monitor_scoreboard_upstream_connection_TB4(1,961,61);
    `monitor_scoreboard_upstream_connection_TB4(1,962,62);
    `monitor_scoreboard_upstream_connection_TB4(1,963,63);
    `monitor_scoreboard_upstream_connection_TB4(1,964,64);
    `monitor_scoreboard_upstream_connection_TB4(1,965,65);
    `monitor_scoreboard_upstream_connection_TB4(1,966,66);
    `monitor_scoreboard_upstream_connection_TB4(1,967,67);
    `monitor_scoreboard_upstream_connection_TB4(1,968,68);
    `monitor_scoreboard_upstream_connection_TB4(1,969,69);
    `monitor_scoreboard_upstream_connection_TB4(1,970,70);
    `monitor_scoreboard_upstream_connection_TB4(1,971,71);
    `monitor_scoreboard_upstream_connection_TB4(1,972,72);
    `monitor_scoreboard_upstream_connection_TB4(1,973,73);
    `monitor_scoreboard_upstream_connection_TB4(1,974,74);
    `monitor_scoreboard_upstream_connection_TB4(1,975,75);
    `monitor_scoreboard_upstream_connection_TB4(1,976,76);
    `monitor_scoreboard_upstream_connection_TB4(1,977,77);
    `monitor_scoreboard_upstream_connection_TB4(1,978,78);
    `monitor_scoreboard_upstream_connection_TB4(1,979,79);
    `monitor_scoreboard_upstream_connection_TB4(1,980,80);
    `monitor_scoreboard_upstream_connection_TB4(1,981,81);
    `monitor_scoreboard_upstream_connection_TB4(1,982,82);
    `monitor_scoreboard_upstream_connection_TB4(1,983,83);
    `monitor_scoreboard_upstream_connection_TB4(1,984,84);
    `monitor_scoreboard_upstream_connection_TB4(1,985,85);
    `monitor_scoreboard_upstream_connection_TB4(1,986,86);
    `monitor_scoreboard_upstream_connection_TB4(1,987,87);
    `monitor_scoreboard_upstream_connection_TB4(1,988,88);
    `monitor_scoreboard_upstream_connection_TB4(1,989,89);
    `monitor_scoreboard_upstream_connection_TB4(1,990,90);
    `monitor_scoreboard_upstream_connection_TB4(1,991,91);
    `monitor_scoreboard_upstream_connection_TB4(1,992,92);
    `monitor_scoreboard_upstream_connection_TB4(1,993,93);
    `monitor_scoreboard_upstream_connection_TB4(1,994,94);
    `monitor_scoreboard_upstream_connection_TB4(1,995,95);
    `monitor_scoreboard_upstream_connection_TB4(1,996,96);
    `monitor_scoreboard_upstream_connection_TB4(1,997,97);
    `monitor_scoreboard_upstream_connection_TB4(1,998,98);
    `monitor_scoreboard_upstream_connection_TB4(1,999,99);
    `monitor_scoreboard_upstream_connection_TB4(1,1000,100);
    `monitor_scoreboard_upstream_connection_TB4(1,1001,101);
    `monitor_scoreboard_upstream_connection_TB4(1,1002,102);
    `monitor_scoreboard_upstream_connection_TB4(1,1003,103);
    `monitor_scoreboard_upstream_connection_TB4(1,1004,104);
    `monitor_scoreboard_upstream_connection_TB4(1,1005,105);
    `monitor_scoreboard_upstream_connection_TB4(1,1006,106);
    `monitor_scoreboard_upstream_connection_TB4(1,1007,107);
    `monitor_scoreboard_upstream_connection_TB4(1,1008,108);
    `monitor_scoreboard_upstream_connection_TB4(1,1009,109);
    `monitor_scoreboard_upstream_connection_TB4(1,1010,110);
    `monitor_scoreboard_upstream_connection_TB4(1,1011,111);
    `monitor_scoreboard_upstream_connection_TB4(1,1012,112);
    `monitor_scoreboard_upstream_connection_TB4(1,1013,113);
    `monitor_scoreboard_upstream_connection_TB4(1,1014,114);
    `monitor_scoreboard_upstream_connection_TB4(1,1015,115);
    `monitor_scoreboard_upstream_connection_TB4(1,1016,116);
    `monitor_scoreboard_upstream_connection_TB4(1,1017,117);
    `monitor_scoreboard_upstream_connection_TB4(1,1018,118);
    `monitor_scoreboard_upstream_connection_TB4(1,1019,119);
    `monitor_scoreboard_upstream_connection_TB4(1,1020,120);
    `monitor_scoreboard_upstream_connection_TB4(1,1021,121);
    `monitor_scoreboard_upstream_connection_TB4(1,1022,122);
    `monitor_scoreboard_upstream_connection_TB4(1,1023,123);
    `monitor_scoreboard_upstream_connection_TB4(1,1024,124);
    `monitor_scoreboard_upstream_connection_TB4(1,1025,125);
    `monitor_scoreboard_upstream_connection_TB4(1,1026,126);
    `monitor_scoreboard_upstream_connection_TB4(1,1027,127);
    `monitor_scoreboard_upstream_connection_TB4(1,1028,128);
    `monitor_scoreboard_upstream_connection_TB4(1,1029,129);
    `monitor_scoreboard_upstream_connection_TB4(1,1030,130);
    `monitor_scoreboard_upstream_connection_TB4(1,1031,131);
    `monitor_scoreboard_upstream_connection_TB4(1,1032,132);
    `monitor_scoreboard_upstream_connection_TB4(1,1033,133);
    `monitor_scoreboard_upstream_connection_TB4(1,1034,134);
    `monitor_scoreboard_upstream_connection_TB4(1,1035,135);
    `monitor_scoreboard_upstream_connection_TB4(1,1036,136);
    `monitor_scoreboard_upstream_connection_TB4(1,1037,137);
    `monitor_scoreboard_upstream_connection_TB4(1,1038,138);
    `monitor_scoreboard_upstream_connection_TB4(1,1039,139);
    `monitor_scoreboard_upstream_connection_TB4(1,1040,140);
    `monitor_scoreboard_upstream_connection_TB4(1,1041,141);
    `monitor_scoreboard_upstream_connection_TB4(1,1042,142);
    `monitor_scoreboard_upstream_connection_TB4(1,1043,143);
    `monitor_scoreboard_upstream_connection_TB4(1,1044,144);
    `monitor_scoreboard_upstream_connection_TB4(1,1045,145);
    `monitor_scoreboard_upstream_connection_TB4(1,1046,146);
    `monitor_scoreboard_upstream_connection_TB4(1,1047,147);
    `monitor_scoreboard_upstream_connection_TB4(1,1048,148);
    `monitor_scoreboard_upstream_connection_TB4(1,1049,149);
    `monitor_scoreboard_upstream_connection_TB4(1,1050,150);
    `monitor_scoreboard_upstream_connection_TB4(1,1051,151);
    `monitor_scoreboard_upstream_connection_TB4(1,1052,152);
    `monitor_scoreboard_upstream_connection_TB4(1,1053,153);
    `monitor_scoreboard_upstream_connection_TB4(1,1054,154);
    `monitor_scoreboard_upstream_connection_TB4(1,1055,155);
    `monitor_scoreboard_upstream_connection_TB4(1,1056,156);
    `monitor_scoreboard_upstream_connection_TB4(1,1057,157);
    `monitor_scoreboard_upstream_connection_TB4(1,1058,158);
    `monitor_scoreboard_upstream_connection_TB4(1,1059,159);
    `monitor_scoreboard_upstream_connection_TB4(1,1060,160);
    `monitor_scoreboard_upstream_connection_TB4(1,1061,161);
    `monitor_scoreboard_upstream_connection_TB4(1,1062,162);
    `monitor_scoreboard_upstream_connection_TB4(1,1063,163);
    `monitor_scoreboard_upstream_connection_TB4(1,1064,164);
    `monitor_scoreboard_upstream_connection_TB4(1,1065,165);
    `monitor_scoreboard_upstream_connection_TB4(1,1066,166);
    `monitor_scoreboard_upstream_connection_TB4(1,1067,167);
    `monitor_scoreboard_upstream_connection_TB4(1,1068,168);
    `monitor_scoreboard_upstream_connection_TB4(1,1069,169);
    `monitor_scoreboard_upstream_connection_TB4(1,1070,170);
    `monitor_scoreboard_upstream_connection_TB4(1,1071,171);
    `monitor_scoreboard_upstream_connection_TB4(1,1072,172);
    `monitor_scoreboard_upstream_connection_TB4(1,1073,173);
    `monitor_scoreboard_upstream_connection_TB4(1,1074,174);
    `monitor_scoreboard_upstream_connection_TB4(1,1075,175);
    `monitor_scoreboard_upstream_connection_TB4(1,1076,176);
    `monitor_scoreboard_upstream_connection_TB4(1,1077,177);
    `monitor_scoreboard_upstream_connection_TB4(1,1078,178);
    `monitor_scoreboard_upstream_connection_TB4(1,1079,179);
    `monitor_scoreboard_upstream_connection_TB4(1,1080,180);
    `monitor_scoreboard_upstream_connection_TB4(1,1081,181);
    `monitor_scoreboard_upstream_connection_TB4(1,1082,182);
    `monitor_scoreboard_upstream_connection_TB4(1,1083,183);
    `monitor_scoreboard_upstream_connection_TB4(1,1084,184);
    `monitor_scoreboard_upstream_connection_TB4(1,1085,185);
    `monitor_scoreboard_upstream_connection_TB4(1,1086,186);
    `monitor_scoreboard_upstream_connection_TB4(1,1087,187);
    `monitor_scoreboard_upstream_connection_TB4(1,1088,188);
    `monitor_scoreboard_upstream_connection_TB4(1,1089,189);
    `monitor_scoreboard_upstream_connection_TB4(1,1090,190);
    `monitor_scoreboard_upstream_connection_TB4(1,1091,191);
    `monitor_scoreboard_upstream_connection_TB4(1,1092,192);
    `monitor_scoreboard_upstream_connection_TB4(1,1093,193);
    `monitor_scoreboard_upstream_connection_TB4(1,1094,194);
    `monitor_scoreboard_upstream_connection_TB4(1,1095,195);
    `monitor_scoreboard_upstream_connection_TB4(1,1096,196);
    `monitor_scoreboard_upstream_connection_TB4(1,1097,197);
    `monitor_scoreboard_upstream_connection_TB4(1,1098,198);
    `monitor_scoreboard_upstream_connection_TB4(1,1099,199);
    `monitor_scoreboard_upstream_connection_TB4(1,1100,200);
    `monitor_scoreboard_upstream_connection_TB4(1,1101,201);
    `monitor_scoreboard_upstream_connection_TB4(1,1102,202);
    `monitor_scoreboard_upstream_connection_TB4(1,1103,203);
    `monitor_scoreboard_upstream_connection_TB4(1,1104,204);
    `monitor_scoreboard_upstream_connection_TB4(1,1105,205);
    `monitor_scoreboard_upstream_connection_TB4(1,1106,206);
    `monitor_scoreboard_upstream_connection_TB4(1,1107,207);
    `monitor_scoreboard_upstream_connection_TB4(1,1108,208);
    `monitor_scoreboard_upstream_connection_TB4(1,1109,209);
    `monitor_scoreboard_upstream_connection_TB4(1,1110,210);
    `monitor_scoreboard_upstream_connection_TB4(1,1111,211);
    `monitor_scoreboard_upstream_connection_TB4(1,1112,212);
    `monitor_scoreboard_upstream_connection_TB4(1,1113,213);
    `monitor_scoreboard_upstream_connection_TB4(1,1114,214);
    `monitor_scoreboard_upstream_connection_TB4(1,1115,215);
    `monitor_scoreboard_upstream_connection_TB4(1,1116,216);
    `monitor_scoreboard_upstream_connection_TB4(1,1117,217);
    `monitor_scoreboard_upstream_connection_TB4(1,1118,218);
    `monitor_scoreboard_upstream_connection_TB4(1,1119,219);
    `monitor_scoreboard_upstream_connection_TB4(1,1120,220);
    `monitor_scoreboard_upstream_connection_TB4(1,1121,221);
    `monitor_scoreboard_upstream_connection_TB4(1,1122,222);
    `monitor_scoreboard_upstream_connection_TB4(1,1123,223);
    `monitor_scoreboard_upstream_connection_TB4(1,1124,224);
    `monitor_scoreboard_upstream_connection_TB4(1,1125,225);
    `monitor_scoreboard_upstream_connection_TB4(1,1126,226);
    `monitor_scoreboard_upstream_connection_TB4(1,1127,227);
    `monitor_scoreboard_upstream_connection_TB4(1,1128,228);
    `monitor_scoreboard_upstream_connection_TB4(1,1129,229);
    `monitor_scoreboard_upstream_connection_TB4(1,1130,230);
    `monitor_scoreboard_upstream_connection_TB4(1,1131,231);
    `monitor_scoreboard_upstream_connection_TB4(1,1132,232);
    `monitor_scoreboard_upstream_connection_TB4(1,1133,233);
    `monitor_scoreboard_upstream_connection_TB4(1,1134,234);
    `monitor_scoreboard_upstream_connection_TB4(1,1135,235);
    `monitor_scoreboard_upstream_connection_TB4(1,1136,236);
    `monitor_scoreboard_upstream_connection_TB4(1,1137,237);
    `monitor_scoreboard_upstream_connection_TB4(1,1138,238);
    `monitor_scoreboard_upstream_connection_TB4(1,1139,239);
    `monitor_scoreboard_upstream_connection_TB4(1,1140,240);
    `monitor_scoreboard_upstream_connection_TB4(1,1141,241);
    `monitor_scoreboard_upstream_connection_TB4(1,1142,242);
    `monitor_scoreboard_upstream_connection_TB4(1,1143,243);
    `monitor_scoreboard_upstream_connection_TB4(1,1144,244);
    `monitor_scoreboard_upstream_connection_TB4(1,1145,245);
    `monitor_scoreboard_upstream_connection_TB4(1,1146,246);
    `monitor_scoreboard_upstream_connection_TB4(1,1147,247);
    `monitor_scoreboard_upstream_connection_TB4(1,1148,248);
    `monitor_scoreboard_upstream_connection_TB4(1,1149,249);
    `monitor_scoreboard_upstream_connection_TB4(1,1150,250);
    `monitor_scoreboard_upstream_connection_TB4(1,1151,251);
    `monitor_scoreboard_upstream_connection_TB4(1,1152,252);
    `monitor_scoreboard_upstream_connection_TB4(1,1153,253);
    `monitor_scoreboard_upstream_connection_TB4(1,1154,254);
    `monitor_scoreboard_upstream_connection_TB4(1,1155,255);
    `monitor_scoreboard_upstream_connection_TB4(1,1156,256);
    `monitor_scoreboard_upstream_connection_TB4(1,1157,257);
    `monitor_scoreboard_upstream_connection_TB4(1,1158,258);
    `monitor_scoreboard_upstream_connection_TB4(1,1159,259);
    `monitor_scoreboard_upstream_connection_TB4(1,1160,260);
    `monitor_scoreboard_upstream_connection_TB4(1,1161,261);
    `monitor_scoreboard_upstream_connection_TB4(1,1162,262);
    `monitor_scoreboard_upstream_connection_TB4(1,1163,263);
    `monitor_scoreboard_upstream_connection_TB4(1,1164,264);
    `monitor_scoreboard_upstream_connection_TB4(1,1165,265);
    `monitor_scoreboard_upstream_connection_TB4(1,1166,266);
    `monitor_scoreboard_upstream_connection_TB4(1,1167,267);
    `monitor_scoreboard_upstream_connection_TB4(1,1168,268);
    `monitor_scoreboard_upstream_connection_TB4(1,1169,269);
    `monitor_scoreboard_upstream_connection_TB4(1,1170,270);
    `monitor_scoreboard_upstream_connection_TB4(1,1171,271);
    `monitor_scoreboard_upstream_connection_TB4(1,1172,272);
    `monitor_scoreboard_upstream_connection_TB4(1,1173,273);
    `monitor_scoreboard_upstream_connection_TB4(1,1174,274);
    `monitor_scoreboard_upstream_connection_TB4(1,1175,275);
    `monitor_scoreboard_upstream_connection_TB4(1,1176,276);
    `monitor_scoreboard_upstream_connection_TB4(1,1177,277);
    `monitor_scoreboard_upstream_connection_TB4(1,1178,278);
    `monitor_scoreboard_upstream_connection_TB4(1,1179,279);
    `monitor_scoreboard_upstream_connection_TB4(1,1180,280);
    `monitor_scoreboard_upstream_connection_TB4(1,1181,281);
    `monitor_scoreboard_upstream_connection_TB4(1,1182,282);
    `monitor_scoreboard_upstream_connection_TB4(1,1183,283);
    `monitor_scoreboard_upstream_connection_TB4(1,1184,284);
    `monitor_scoreboard_upstream_connection_TB4(1,1185,285);
    `monitor_scoreboard_upstream_connection_TB4(1,1186,286);
    `monitor_scoreboard_upstream_connection_TB4(1,1187,287);
    `monitor_scoreboard_upstream_connection_TB4(1,1188,288);
    `monitor_scoreboard_upstream_connection_TB4(1,1189,289);
    `monitor_scoreboard_upstream_connection_TB4(1,1190,290);
    `monitor_scoreboard_upstream_connection_TB4(1,1191,291);
    `monitor_scoreboard_upstream_connection_TB4(1,1192,292);
    `monitor_scoreboard_upstream_connection_TB4(1,1193,293);
    `monitor_scoreboard_upstream_connection_TB4(1,1194,294);
    `monitor_scoreboard_upstream_connection_TB4(1,1195,295);
    `monitor_scoreboard_upstream_connection_TB4(1,1196,296);
    `monitor_scoreboard_upstream_connection_TB4(1,1197,297);
    `monitor_scoreboard_upstream_connection_TB4(1,1198,298);
    `monitor_scoreboard_upstream_connection_TB4(1,1199,299);
    `monitor_scoreboard_upstream_connection_TB4(1,1200,300);
    `monitor_scoreboard_upstream_connection_TB4(1,1201,301);
    `monitor_scoreboard_upstream_connection_TB4(1,1202,302);
    `monitor_scoreboard_upstream_connection_TB4(1,1203,303);
    `monitor_scoreboard_upstream_connection_TB4(1,1204,304);
    `monitor_scoreboard_upstream_connection_TB4(1,1205,305);
    `monitor_scoreboard_upstream_connection_TB4(1,1206,306);
    `monitor_scoreboard_upstream_connection_TB4(1,1207,307);
    `monitor_scoreboard_upstream_connection_TB4(1,1208,308);
    `monitor_scoreboard_upstream_connection_TB4(1,1209,309);
    `monitor_scoreboard_upstream_connection_TB4(1,1210,310);
    `monitor_scoreboard_upstream_connection_TB4(1,1211,311);
    `monitor_scoreboard_upstream_connection_TB4(1,1212,312);
    `monitor_scoreboard_upstream_connection_TB4(1,1213,313);
    `monitor_scoreboard_upstream_connection_TB4(1,1214,314);
    `monitor_scoreboard_upstream_connection_TB4(1,1215,315);
    `monitor_scoreboard_upstream_connection_TB4(1,1216,316);
    `monitor_scoreboard_upstream_connection_TB4(1,1217,317);
    `monitor_scoreboard_upstream_connection_TB4(1,1218,318);
    `monitor_scoreboard_upstream_connection_TB4(1,1219,319);
    `monitor_scoreboard_upstream_connection_TB4(1,1220,320);
    `monitor_scoreboard_upstream_connection_TB4(1,1221,321);
    `monitor_scoreboard_upstream_connection_TB4(1,1222,322);
    `monitor_scoreboard_upstream_connection_TB4(1,1223,323);
    `monitor_scoreboard_upstream_connection_TB4(1,1224,324);
    `monitor_scoreboard_upstream_connection_TB4(1,1225,325);
    `monitor_scoreboard_upstream_connection_TB4(1,1226,326);
    `monitor_scoreboard_upstream_connection_TB4(1,1227,327);
    `monitor_scoreboard_upstream_connection_TB4(1,1228,328);
    `monitor_scoreboard_upstream_connection_TB4(1,1229,329);
    `monitor_scoreboard_upstream_connection_TB4(1,1230,330);
    `monitor_scoreboard_upstream_connection_TB4(1,1231,331);
    `monitor_scoreboard_upstream_connection_TB4(1,1232,332);
    `monitor_scoreboard_upstream_connection_TB4(1,1233,333);
    `monitor_scoreboard_upstream_connection_TB4(1,1234,334);
    `monitor_scoreboard_upstream_connection_TB4(1,1235,335);
    `monitor_scoreboard_upstream_connection_TB4(1,1236,336);
    `monitor_scoreboard_upstream_connection_TB4(1,1237,337);
    `monitor_scoreboard_upstream_connection_TB4(1,1238,338);
    `monitor_scoreboard_upstream_connection_TB4(1,1239,339);
    `monitor_scoreboard_upstream_connection_TB4(1,1240,340);
    `monitor_scoreboard_upstream_connection_TB4(1,1241,341);
    `monitor_scoreboard_upstream_connection_TB4(1,1242,342);
    `monitor_scoreboard_upstream_connection_TB4(1,1243,343);
    `monitor_scoreboard_upstream_connection_TB4(1,1244,344);
    `monitor_scoreboard_upstream_connection_TB4(1,1245,345);
    `monitor_scoreboard_upstream_connection_TB4(1,1246,346);
    `monitor_scoreboard_upstream_connection_TB4(1,1247,347);
    `monitor_scoreboard_upstream_connection_TB4(1,1248,348);
    `monitor_scoreboard_upstream_connection_TB4(1,1249,349);
    `monitor_scoreboard_upstream_connection_TB4(1,1250,350);
    `monitor_scoreboard_upstream_connection_TB4(1,1251,351);
    `monitor_scoreboard_upstream_connection_TB4(1,1252,352);
    `monitor_scoreboard_upstream_connection_TB4(1,1253,353);
    `monitor_scoreboard_upstream_connection_TB4(1,1254,354);
    `monitor_scoreboard_upstream_connection_TB4(1,1255,355);
    `monitor_scoreboard_upstream_connection_TB4(1,1256,356);
    `monitor_scoreboard_upstream_connection_TB4(1,1257,357);
    `monitor_scoreboard_upstream_connection_TB4(1,1258,358);
    `monitor_scoreboard_upstream_connection_TB4(1,1259,359);
    `monitor_scoreboard_upstream_connection_TB4(1,1260,360);
    `monitor_scoreboard_upstream_connection_TB4(1,1261,361);
    `monitor_scoreboard_upstream_connection_TB4(1,1262,362);
    `monitor_scoreboard_upstream_connection_TB4(1,1263,363);
    `monitor_scoreboard_upstream_connection_TB4(1,1264,364);
    `monitor_scoreboard_upstream_connection_TB4(1,1265,365);
    `monitor_scoreboard_upstream_connection_TB4(1,1266,366);
    `monitor_scoreboard_upstream_connection_TB4(1,1267,367);
    `monitor_scoreboard_upstream_connection_TB4(1,1268,368);
    `monitor_scoreboard_upstream_connection_TB4(1,1269,369);
    `monitor_scoreboard_upstream_connection_TB4(1,1270,370);
    `monitor_scoreboard_upstream_connection_TB4(1,1271,371);
    `monitor_scoreboard_upstream_connection_TB4(1,1272,372);
    `monitor_scoreboard_upstream_connection_TB4(1,1273,373);
    `monitor_scoreboard_upstream_connection_TB4(1,1274,374);
    `monitor_scoreboard_upstream_connection_TB4(1,1275,375);
    `monitor_scoreboard_upstream_connection_TB4(1,1276,376);
    `monitor_scoreboard_upstream_connection_TB4(1,1277,377);
    `monitor_scoreboard_upstream_connection_TB4(1,1278,378);
    `monitor_scoreboard_upstream_connection_TB4(1,1279,379);
    `monitor_scoreboard_upstream_connection_TB4(1,1280,380);
    `monitor_scoreboard_upstream_connection_TB4(1,1281,381);
    `monitor_scoreboard_upstream_connection_TB4(1,1282,382);
    `monitor_scoreboard_upstream_connection_TB4(1,1283,383);
    `monitor_scoreboard_upstream_connection_TB4(1,1284,384);
    `monitor_scoreboard_upstream_connection_TB4(1,1285,385);
    `monitor_scoreboard_upstream_connection_TB4(1,1286,386);
    `monitor_scoreboard_upstream_connection_TB4(1,1287,387);
    `monitor_scoreboard_upstream_connection_TB4(1,1288,388);
    `monitor_scoreboard_upstream_connection_TB4(1,1289,389);
    `monitor_scoreboard_upstream_connection_TB4(1,1290,390);
    `monitor_scoreboard_upstream_connection_TB4(1,1291,391);
    `monitor_scoreboard_upstream_connection_TB4(1,1292,392);
    `monitor_scoreboard_upstream_connection_TB4(1,1293,393);
    `monitor_scoreboard_upstream_connection_TB4(1,1294,394);
    `monitor_scoreboard_upstream_connection_TB4(1,1295,395);
    `monitor_scoreboard_upstream_connection_TB4(1,1296,396);
    `monitor_scoreboard_upstream_connection_TB4(1,1297,397);
    `monitor_scoreboard_upstream_connection_TB4(1,1298,398);
    `monitor_scoreboard_upstream_connection_TB4(1,1299,399);
    `monitor_scoreboard_upstream_connection_TB4(1,1300,400);
    `monitor_scoreboard_upstream_connection_TB4(1,1301,401);
    `monitor_scoreboard_upstream_connection_TB4(1,1302,402);
    `monitor_scoreboard_upstream_connection_TB4(1,1303,403);
    `monitor_scoreboard_upstream_connection_TB4(1,1304,404);
    `monitor_scoreboard_upstream_connection_TB4(1,1305,405);
    `monitor_scoreboard_upstream_connection_TB4(1,1306,406);
    `monitor_scoreboard_upstream_connection_TB4(1,1307,407);
    `monitor_scoreboard_upstream_connection_TB4(1,1308,408);
    `monitor_scoreboard_upstream_connection_TB4(1,1309,409);
    `monitor_scoreboard_upstream_connection_TB4(1,1310,410);
    `monitor_scoreboard_upstream_connection_TB4(1,1311,411);
    `monitor_scoreboard_upstream_connection_TB4(1,1312,412);
    `monitor_scoreboard_upstream_connection_TB4(1,1313,413);
    `monitor_scoreboard_upstream_connection_TB4(1,1314,414);
    `monitor_scoreboard_upstream_connection_TB4(1,1315,415);
    `monitor_scoreboard_upstream_connection_TB4(1,1316,416);
    `monitor_scoreboard_upstream_connection_TB4(1,1317,417);
    `monitor_scoreboard_upstream_connection_TB4(1,1318,418);
    `monitor_scoreboard_upstream_connection_TB4(1,1319,419);
    `monitor_scoreboard_upstream_connection_TB4(1,1320,420);
    `monitor_scoreboard_upstream_connection_TB4(1,1321,421);
    `monitor_scoreboard_upstream_connection_TB4(1,1322,422);
    `monitor_scoreboard_upstream_connection_TB4(1,1323,423);
    `monitor_scoreboard_upstream_connection_TB4(1,1324,424);
    `monitor_scoreboard_upstream_connection_TB4(1,1325,425);
    `monitor_scoreboard_upstream_connection_TB4(1,1326,426);
    `monitor_scoreboard_upstream_connection_TB4(1,1327,427);
    `monitor_scoreboard_upstream_connection_TB4(1,1328,428);
    `monitor_scoreboard_upstream_connection_TB4(1,1329,429);
    `monitor_scoreboard_upstream_connection_TB4(1,1330,430);
    `monitor_scoreboard_upstream_connection_TB4(1,1331,431);
    `monitor_scoreboard_upstream_connection_TB4(1,1332,432);
    `monitor_scoreboard_upstream_connection_TB4(1,1333,433);
    `monitor_scoreboard_upstream_connection_TB4(1,1334,434);
    `monitor_scoreboard_upstream_connection_TB4(1,1335,435);
    `monitor_scoreboard_upstream_connection_TB4(1,1336,436);
    `monitor_scoreboard_upstream_connection_TB4(1,1337,437);
    `monitor_scoreboard_upstream_connection_TB4(1,1338,438);
    `monitor_scoreboard_upstream_connection_TB4(1,1339,439);
    `monitor_scoreboard_upstream_connection_TB4(1,1340,440);
    `monitor_scoreboard_upstream_connection_TB4(1,1341,441);
    `monitor_scoreboard_upstream_connection_TB4(1,1342,442);
    `monitor_scoreboard_upstream_connection_TB4(1,1343,443);
    `monitor_scoreboard_upstream_connection_TB4(1,1344,444);
    `monitor_scoreboard_upstream_connection_TB4(1,1345,445);
    `monitor_scoreboard_upstream_connection_TB4(1,1346,446);
    `monitor_scoreboard_upstream_connection_TB4(1,1347,447);
    `monitor_scoreboard_upstream_connection_TB4(1,1348,448);
    `monitor_scoreboard_upstream_connection_TB4(1,1349,449);
    `monitor_scoreboard_upstream_connection_TB4(2,1350,0);
    `monitor_scoreboard_upstream_connection_TB4(2,1351,1);
    `monitor_scoreboard_upstream_connection_TB4(2,1352,2);
    `monitor_scoreboard_upstream_connection_TB4(2,1353,3);
    `monitor_scoreboard_upstream_connection_TB4(2,1354,4);
    `monitor_scoreboard_upstream_connection_TB4(2,1355,5);
    `monitor_scoreboard_upstream_connection_TB4(2,1356,6);
    `monitor_scoreboard_upstream_connection_TB4(2,1357,7);
    `monitor_scoreboard_upstream_connection_TB4(2,1358,8);
    `monitor_scoreboard_upstream_connection_TB4(2,1359,9);
    `monitor_scoreboard_upstream_connection_TB4(2,1360,10);
    `monitor_scoreboard_upstream_connection_TB4(2,1361,11);
    `monitor_scoreboard_upstream_connection_TB4(2,1362,12);
    `monitor_scoreboard_upstream_connection_TB4(2,1363,13);
    `monitor_scoreboard_upstream_connection_TB4(2,1364,14);
    `monitor_scoreboard_upstream_connection_TB4(2,1365,15);
    `monitor_scoreboard_upstream_connection_TB4(2,1366,16);
    `monitor_scoreboard_upstream_connection_TB4(2,1367,17);
    `monitor_scoreboard_upstream_connection_TB4(2,1368,18);
    `monitor_scoreboard_upstream_connection_TB4(2,1369,19);
    `monitor_scoreboard_upstream_connection_TB4(2,1370,20);
    `monitor_scoreboard_upstream_connection_TB4(2,1371,21);
    `monitor_scoreboard_upstream_connection_TB4(2,1372,22);
    `monitor_scoreboard_upstream_connection_TB4(2,1373,23);
    `monitor_scoreboard_upstream_connection_TB4(2,1374,24);
    `monitor_scoreboard_upstream_connection_TB4(2,1375,25);
    `monitor_scoreboard_upstream_connection_TB4(2,1376,26);
    `monitor_scoreboard_upstream_connection_TB4(2,1377,27);
    `monitor_scoreboard_upstream_connection_TB4(2,1378,28);
    `monitor_scoreboard_upstream_connection_TB4(2,1379,29);
    `monitor_scoreboard_upstream_connection_TB4(2,1380,30);
    `monitor_scoreboard_upstream_connection_TB4(2,1381,31);
    `monitor_scoreboard_upstream_connection_TB4(2,1382,32);
    `monitor_scoreboard_upstream_connection_TB4(2,1383,33);
    `monitor_scoreboard_upstream_connection_TB4(2,1384,34);
    `monitor_scoreboard_upstream_connection_TB4(2,1385,35);
    `monitor_scoreboard_upstream_connection_TB4(2,1386,36);
    `monitor_scoreboard_upstream_connection_TB4(2,1387,37);
    `monitor_scoreboard_upstream_connection_TB4(2,1388,38);
    `monitor_scoreboard_upstream_connection_TB4(2,1389,39);
    `monitor_scoreboard_upstream_connection_TB4(2,1390,40);
    `monitor_scoreboard_upstream_connection_TB4(2,1391,41);
    `monitor_scoreboard_upstream_connection_TB4(2,1392,42);
    `monitor_scoreboard_upstream_connection_TB4(2,1393,43);
    `monitor_scoreboard_upstream_connection_TB4(2,1394,44);
    `monitor_scoreboard_upstream_connection_TB4(2,1395,45);
    `monitor_scoreboard_upstream_connection_TB4(2,1396,46);
    `monitor_scoreboard_upstream_connection_TB4(2,1397,47);
    `monitor_scoreboard_upstream_connection_TB4(2,1398,48);
    `monitor_scoreboard_upstream_connection_TB4(2,1399,49);
    `monitor_scoreboard_upstream_connection_TB4(2,1400,50);
    `monitor_scoreboard_upstream_connection_TB4(2,1401,51);
    `monitor_scoreboard_upstream_connection_TB4(2,1402,52);
    `monitor_scoreboard_upstream_connection_TB4(2,1403,53);
    `monitor_scoreboard_upstream_connection_TB4(2,1404,54);
    `monitor_scoreboard_upstream_connection_TB4(2,1405,55);
    `monitor_scoreboard_upstream_connection_TB4(2,1406,56);
    `monitor_scoreboard_upstream_connection_TB4(2,1407,57);
    `monitor_scoreboard_upstream_connection_TB4(2,1408,58);
    `monitor_scoreboard_upstream_connection_TB4(2,1409,59);
    `monitor_scoreboard_upstream_connection_TB4(2,1410,60);
    `monitor_scoreboard_upstream_connection_TB4(2,1411,61);
    `monitor_scoreboard_upstream_connection_TB4(2,1412,62);
    `monitor_scoreboard_upstream_connection_TB4(2,1413,63);
    `monitor_scoreboard_upstream_connection_TB4(2,1414,64);
    `monitor_scoreboard_upstream_connection_TB4(2,1415,65);
    `monitor_scoreboard_upstream_connection_TB4(2,1416,66);
    `monitor_scoreboard_upstream_connection_TB4(2,1417,67);
    `monitor_scoreboard_upstream_connection_TB4(2,1418,68);
    `monitor_scoreboard_upstream_connection_TB4(2,1419,69);
    `monitor_scoreboard_upstream_connection_TB4(2,1420,70);
    `monitor_scoreboard_upstream_connection_TB4(2,1421,71);
    `monitor_scoreboard_upstream_connection_TB4(2,1422,72);
    `monitor_scoreboard_upstream_connection_TB4(2,1423,73);
    `monitor_scoreboard_upstream_connection_TB4(2,1424,74);
    `monitor_scoreboard_upstream_connection_TB4(2,1425,75);
    `monitor_scoreboard_upstream_connection_TB4(2,1426,76);
    `monitor_scoreboard_upstream_connection_TB4(2,1427,77);
    `monitor_scoreboard_upstream_connection_TB4(2,1428,78);
    `monitor_scoreboard_upstream_connection_TB4(2,1429,79);
    `monitor_scoreboard_upstream_connection_TB4(2,1430,80);
    `monitor_scoreboard_upstream_connection_TB4(2,1431,81);
    `monitor_scoreboard_upstream_connection_TB4(2,1432,82);
    `monitor_scoreboard_upstream_connection_TB4(2,1433,83);
    `monitor_scoreboard_upstream_connection_TB4(2,1434,84);
    `monitor_scoreboard_upstream_connection_TB4(2,1435,85);
    `monitor_scoreboard_upstream_connection_TB4(2,1436,86);
    `monitor_scoreboard_upstream_connection_TB4(2,1437,87);
    `monitor_scoreboard_upstream_connection_TB4(2,1438,88);
    `monitor_scoreboard_upstream_connection_TB4(2,1439,89);
    `monitor_scoreboard_upstream_connection_TB4(2,1440,90);
    `monitor_scoreboard_upstream_connection_TB4(2,1441,91);
    `monitor_scoreboard_upstream_connection_TB4(2,1442,92);
    `monitor_scoreboard_upstream_connection_TB4(2,1443,93);
    `monitor_scoreboard_upstream_connection_TB4(2,1444,94);
    `monitor_scoreboard_upstream_connection_TB4(2,1445,95);
    `monitor_scoreboard_upstream_connection_TB4(2,1446,96);
    `monitor_scoreboard_upstream_connection_TB4(2,1447,97);
    `monitor_scoreboard_upstream_connection_TB4(2,1448,98);
    `monitor_scoreboard_upstream_connection_TB4(2,1449,99);
    `monitor_scoreboard_upstream_connection_TB4(2,1450,100);
    `monitor_scoreboard_upstream_connection_TB4(2,1451,101);
    `monitor_scoreboard_upstream_connection_TB4(2,1452,102);
    `monitor_scoreboard_upstream_connection_TB4(2,1453,103);
    `monitor_scoreboard_upstream_connection_TB4(2,1454,104);
    `monitor_scoreboard_upstream_connection_TB4(2,1455,105);
    `monitor_scoreboard_upstream_connection_TB4(2,1456,106);
    `monitor_scoreboard_upstream_connection_TB4(2,1457,107);
    `monitor_scoreboard_upstream_connection_TB4(2,1458,108);
    `monitor_scoreboard_upstream_connection_TB4(2,1459,109);
    `monitor_scoreboard_upstream_connection_TB4(2,1460,110);
    `monitor_scoreboard_upstream_connection_TB4(2,1461,111);
    `monitor_scoreboard_upstream_connection_TB4(2,1462,112);
    `monitor_scoreboard_upstream_connection_TB4(2,1463,113);
    `monitor_scoreboard_upstream_connection_TB4(2,1464,114);
    `monitor_scoreboard_upstream_connection_TB4(2,1465,115);
    `monitor_scoreboard_upstream_connection_TB4(2,1466,116);
    `monitor_scoreboard_upstream_connection_TB4(2,1467,117);
    `monitor_scoreboard_upstream_connection_TB4(2,1468,118);
    `monitor_scoreboard_upstream_connection_TB4(2,1469,119);
    `monitor_scoreboard_upstream_connection_TB4(2,1470,120);
    `monitor_scoreboard_upstream_connection_TB4(2,1471,121);
    `monitor_scoreboard_upstream_connection_TB4(2,1472,122);
    `monitor_scoreboard_upstream_connection_TB4(2,1473,123);
    `monitor_scoreboard_upstream_connection_TB4(2,1474,124);
    `monitor_scoreboard_upstream_connection_TB4(2,1475,125);
    `monitor_scoreboard_upstream_connection_TB4(2,1476,126);
    `monitor_scoreboard_upstream_connection_TB4(2,1477,127);
    `monitor_scoreboard_upstream_connection_TB4(2,1478,128);
    `monitor_scoreboard_upstream_connection_TB4(2,1479,129);
    `monitor_scoreboard_upstream_connection_TB4(2,1480,130);
    `monitor_scoreboard_upstream_connection_TB4(2,1481,131);
    `monitor_scoreboard_upstream_connection_TB4(2,1482,132);
    `monitor_scoreboard_upstream_connection_TB4(2,1483,133);
    `monitor_scoreboard_upstream_connection_TB4(2,1484,134);
    `monitor_scoreboard_upstream_connection_TB4(2,1485,135);
    `monitor_scoreboard_upstream_connection_TB4(2,1486,136);
    `monitor_scoreboard_upstream_connection_TB4(2,1487,137);
    `monitor_scoreboard_upstream_connection_TB4(2,1488,138);
    `monitor_scoreboard_upstream_connection_TB4(2,1489,139);
    `monitor_scoreboard_upstream_connection_TB4(2,1490,140);
    `monitor_scoreboard_upstream_connection_TB4(2,1491,141);
    `monitor_scoreboard_upstream_connection_TB4(2,1492,142);
    `monitor_scoreboard_upstream_connection_TB4(2,1493,143);
    `monitor_scoreboard_upstream_connection_TB4(2,1494,144);
    `monitor_scoreboard_upstream_connection_TB4(2,1495,145);
    `monitor_scoreboard_upstream_connection_TB4(2,1496,146);
    `monitor_scoreboard_upstream_connection_TB4(2,1497,147);
    `monitor_scoreboard_upstream_connection_TB4(2,1498,148);
    `monitor_scoreboard_upstream_connection_TB4(2,1499,149);
    `monitor_scoreboard_upstream_connection_TB4(2,1500,150);
    `monitor_scoreboard_upstream_connection_TB4(2,1501,151);
    `monitor_scoreboard_upstream_connection_TB4(2,1502,152);
    `monitor_scoreboard_upstream_connection_TB4(2,1503,153);
    `monitor_scoreboard_upstream_connection_TB4(2,1504,154);
    `monitor_scoreboard_upstream_connection_TB4(2,1505,155);
    `monitor_scoreboard_upstream_connection_TB4(2,1506,156);
    `monitor_scoreboard_upstream_connection_TB4(2,1507,157);
    `monitor_scoreboard_upstream_connection_TB4(2,1508,158);
    `monitor_scoreboard_upstream_connection_TB4(2,1509,159);
    `monitor_scoreboard_upstream_connection_TB4(2,1510,160);
    `monitor_scoreboard_upstream_connection_TB4(2,1511,161);
    `monitor_scoreboard_upstream_connection_TB4(2,1512,162);
    `monitor_scoreboard_upstream_connection_TB4(2,1513,163);
    `monitor_scoreboard_upstream_connection_TB4(2,1514,164);
    `monitor_scoreboard_upstream_connection_TB4(2,1515,165);
    `monitor_scoreboard_upstream_connection_TB4(2,1516,166);
    `monitor_scoreboard_upstream_connection_TB4(2,1517,167);
    `monitor_scoreboard_upstream_connection_TB4(2,1518,168);
    `monitor_scoreboard_upstream_connection_TB4(2,1519,169);
    `monitor_scoreboard_upstream_connection_TB4(2,1520,170);
    `monitor_scoreboard_upstream_connection_TB4(2,1521,171);
    `monitor_scoreboard_upstream_connection_TB4(2,1522,172);
    `monitor_scoreboard_upstream_connection_TB4(2,1523,173);
    `monitor_scoreboard_upstream_connection_TB4(2,1524,174);
    `monitor_scoreboard_upstream_connection_TB4(2,1525,175);
    `monitor_scoreboard_upstream_connection_TB4(2,1526,176);
    `monitor_scoreboard_upstream_connection_TB4(2,1527,177);
    `monitor_scoreboard_upstream_connection_TB4(2,1528,178);
    `monitor_scoreboard_upstream_connection_TB4(2,1529,179);
    `monitor_scoreboard_upstream_connection_TB4(2,1530,180);
    `monitor_scoreboard_upstream_connection_TB4(2,1531,181);
    `monitor_scoreboard_upstream_connection_TB4(2,1532,182);
    `monitor_scoreboard_upstream_connection_TB4(2,1533,183);
    `monitor_scoreboard_upstream_connection_TB4(2,1534,184);
    `monitor_scoreboard_upstream_connection_TB4(2,1535,185);
    `monitor_scoreboard_upstream_connection_TB4(2,1536,186);
    `monitor_scoreboard_upstream_connection_TB4(2,1537,187);
    `monitor_scoreboard_upstream_connection_TB4(2,1538,188);
    `monitor_scoreboard_upstream_connection_TB4(2,1539,189);
    `monitor_scoreboard_upstream_connection_TB4(2,1540,190);
    `monitor_scoreboard_upstream_connection_TB4(2,1541,191);
    `monitor_scoreboard_upstream_connection_TB4(2,1542,192);
    `monitor_scoreboard_upstream_connection_TB4(2,1543,193);
    `monitor_scoreboard_upstream_connection_TB4(2,1544,194);
    `monitor_scoreboard_upstream_connection_TB4(2,1545,195);
    `monitor_scoreboard_upstream_connection_TB4(2,1546,196);
    `monitor_scoreboard_upstream_connection_TB4(2,1547,197);
    `monitor_scoreboard_upstream_connection_TB4(2,1548,198);
    `monitor_scoreboard_upstream_connection_TB4(2,1549,199);
    `monitor_scoreboard_upstream_connection_TB4(2,1550,200);
    `monitor_scoreboard_upstream_connection_TB4(2,1551,201);
    `monitor_scoreboard_upstream_connection_TB4(2,1552,202);
    `monitor_scoreboard_upstream_connection_TB4(2,1553,203);
    `monitor_scoreboard_upstream_connection_TB4(2,1554,204);
    `monitor_scoreboard_upstream_connection_TB4(2,1555,205);
    `monitor_scoreboard_upstream_connection_TB4(2,1556,206);
    `monitor_scoreboard_upstream_connection_TB4(2,1557,207);
    `monitor_scoreboard_upstream_connection_TB4(2,1558,208);
    `monitor_scoreboard_upstream_connection_TB4(2,1559,209);
    `monitor_scoreboard_upstream_connection_TB4(2,1560,210);
    `monitor_scoreboard_upstream_connection_TB4(2,1561,211);
    `monitor_scoreboard_upstream_connection_TB4(2,1562,212);
    `monitor_scoreboard_upstream_connection_TB4(2,1563,213);
    `monitor_scoreboard_upstream_connection_TB4(2,1564,214);
    `monitor_scoreboard_upstream_connection_TB4(2,1565,215);
    `monitor_scoreboard_upstream_connection_TB4(2,1566,216);
    `monitor_scoreboard_upstream_connection_TB4(2,1567,217);
    `monitor_scoreboard_upstream_connection_TB4(2,1568,218);
    `monitor_scoreboard_upstream_connection_TB4(2,1569,219);
    `monitor_scoreboard_upstream_connection_TB4(2,1570,220);
    `monitor_scoreboard_upstream_connection_TB4(2,1571,221);
    `monitor_scoreboard_upstream_connection_TB4(2,1572,222);
    `monitor_scoreboard_upstream_connection_TB4(2,1573,223);
    `monitor_scoreboard_upstream_connection_TB4(2,1574,224);
    `monitor_scoreboard_upstream_connection_TB4(2,1575,225);
    `monitor_scoreboard_upstream_connection_TB4(2,1576,226);
    `monitor_scoreboard_upstream_connection_TB4(2,1577,227);
    `monitor_scoreboard_upstream_connection_TB4(2,1578,228);
    `monitor_scoreboard_upstream_connection_TB4(2,1579,229);
    `monitor_scoreboard_upstream_connection_TB4(2,1580,230);
    `monitor_scoreboard_upstream_connection_TB4(2,1581,231);
    `monitor_scoreboard_upstream_connection_TB4(2,1582,232);
    `monitor_scoreboard_upstream_connection_TB4(2,1583,233);
    `monitor_scoreboard_upstream_connection_TB4(2,1584,234);
    `monitor_scoreboard_upstream_connection_TB4(2,1585,235);
    `monitor_scoreboard_upstream_connection_TB4(2,1586,236);
    `monitor_scoreboard_upstream_connection_TB4(2,1587,237);
    `monitor_scoreboard_upstream_connection_TB4(2,1588,238);
    `monitor_scoreboard_upstream_connection_TB4(2,1589,239);
    `monitor_scoreboard_upstream_connection_TB4(2,1590,240);
    `monitor_scoreboard_upstream_connection_TB4(2,1591,241);
    `monitor_scoreboard_upstream_connection_TB4(2,1592,242);
    `monitor_scoreboard_upstream_connection_TB4(2,1593,243);
    `monitor_scoreboard_upstream_connection_TB4(2,1594,244);
    `monitor_scoreboard_upstream_connection_TB4(2,1595,245);
    `monitor_scoreboard_upstream_connection_TB4(2,1596,246);
    `monitor_scoreboard_upstream_connection_TB4(2,1597,247);
    `monitor_scoreboard_upstream_connection_TB4(2,1598,248);
    `monitor_scoreboard_upstream_connection_TB4(2,1599,249);
    `monitor_scoreboard_upstream_connection_TB4(2,1600,250);
    `monitor_scoreboard_upstream_connection_TB4(2,1601,251);
    `monitor_scoreboard_upstream_connection_TB4(2,1602,252);
    `monitor_scoreboard_upstream_connection_TB4(2,1603,253);
    `monitor_scoreboard_upstream_connection_TB4(2,1604,254);
    `monitor_scoreboard_upstream_connection_TB4(2,1605,255);
    `monitor_scoreboard_upstream_connection_TB4(2,1606,256);
    `monitor_scoreboard_upstream_connection_TB4(2,1607,257);
    `monitor_scoreboard_upstream_connection_TB4(2,1608,258);
    `monitor_scoreboard_upstream_connection_TB4(2,1609,259);
    `monitor_scoreboard_upstream_connection_TB4(2,1610,260);
    `monitor_scoreboard_upstream_connection_TB4(2,1611,261);
    `monitor_scoreboard_upstream_connection_TB4(2,1612,262);
    `monitor_scoreboard_upstream_connection_TB4(2,1613,263);
    `monitor_scoreboard_upstream_connection_TB4(2,1614,264);
    `monitor_scoreboard_upstream_connection_TB4(2,1615,265);
    `monitor_scoreboard_upstream_connection_TB4(2,1616,266);
    `monitor_scoreboard_upstream_connection_TB4(2,1617,267);
    `monitor_scoreboard_upstream_connection_TB4(2,1618,268);
    `monitor_scoreboard_upstream_connection_TB4(2,1619,269);
    `monitor_scoreboard_upstream_connection_TB4(2,1620,270);
    `monitor_scoreboard_upstream_connection_TB4(2,1621,271);
    `monitor_scoreboard_upstream_connection_TB4(2,1622,272);
    `monitor_scoreboard_upstream_connection_TB4(2,1623,273);
    `monitor_scoreboard_upstream_connection_TB4(2,1624,274);
    `monitor_scoreboard_upstream_connection_TB4(2,1625,275);
    `monitor_scoreboard_upstream_connection_TB4(2,1626,276);
    `monitor_scoreboard_upstream_connection_TB4(2,1627,277);
    `monitor_scoreboard_upstream_connection_TB4(2,1628,278);
    `monitor_scoreboard_upstream_connection_TB4(2,1629,279);
    `monitor_scoreboard_upstream_connection_TB4(2,1630,280);
    `monitor_scoreboard_upstream_connection_TB4(2,1631,281);
    `monitor_scoreboard_upstream_connection_TB4(2,1632,282);
    `monitor_scoreboard_upstream_connection_TB4(2,1633,283);
    `monitor_scoreboard_upstream_connection_TB4(2,1634,284);
    `monitor_scoreboard_upstream_connection_TB4(2,1635,285);
    `monitor_scoreboard_upstream_connection_TB4(2,1636,286);
    `monitor_scoreboard_upstream_connection_TB4(2,1637,287);
    `monitor_scoreboard_upstream_connection_TB4(2,1638,288);
    `monitor_scoreboard_upstream_connection_TB4(2,1639,289);
    `monitor_scoreboard_upstream_connection_TB4(2,1640,290);
    `monitor_scoreboard_upstream_connection_TB4(2,1641,291);
    `monitor_scoreboard_upstream_connection_TB4(2,1642,292);
    `monitor_scoreboard_upstream_connection_TB4(2,1643,293);
    `monitor_scoreboard_upstream_connection_TB4(2,1644,294);
    `monitor_scoreboard_upstream_connection_TB4(2,1645,295);
    `monitor_scoreboard_upstream_connection_TB4(2,1646,296);
    `monitor_scoreboard_upstream_connection_TB4(2,1647,297);
    `monitor_scoreboard_upstream_connection_TB4(2,1648,298);
    `monitor_scoreboard_upstream_connection_TB4(2,1649,299);
    `monitor_scoreboard_upstream_connection_TB4(2,1650,300);
    `monitor_scoreboard_upstream_connection_TB4(2,1651,301);
    `monitor_scoreboard_upstream_connection_TB4(2,1652,302);
    `monitor_scoreboard_upstream_connection_TB4(2,1653,303);
    `monitor_scoreboard_upstream_connection_TB4(2,1654,304);
    `monitor_scoreboard_upstream_connection_TB4(2,1655,305);
    `monitor_scoreboard_upstream_connection_TB4(2,1656,306);
    `monitor_scoreboard_upstream_connection_TB4(2,1657,307);
    `monitor_scoreboard_upstream_connection_TB4(2,1658,308);
    `monitor_scoreboard_upstream_connection_TB4(2,1659,309);
    `monitor_scoreboard_upstream_connection_TB4(2,1660,310);
    `monitor_scoreboard_upstream_connection_TB4(2,1661,311);
    `monitor_scoreboard_upstream_connection_TB4(2,1662,312);
    `monitor_scoreboard_upstream_connection_TB4(2,1663,313);
    `monitor_scoreboard_upstream_connection_TB4(2,1664,314);
    `monitor_scoreboard_upstream_connection_TB4(2,1665,315);
    `monitor_scoreboard_upstream_connection_TB4(2,1666,316);
    `monitor_scoreboard_upstream_connection_TB4(2,1667,317);
    `monitor_scoreboard_upstream_connection_TB4(2,1668,318);
    `monitor_scoreboard_upstream_connection_TB4(2,1669,319);
    `monitor_scoreboard_upstream_connection_TB4(2,1670,320);
    `monitor_scoreboard_upstream_connection_TB4(2,1671,321);
    `monitor_scoreboard_upstream_connection_TB4(2,1672,322);
    `monitor_scoreboard_upstream_connection_TB4(2,1673,323);
    `monitor_scoreboard_upstream_connection_TB4(2,1674,324);
    `monitor_scoreboard_upstream_connection_TB4(2,1675,325);
    `monitor_scoreboard_upstream_connection_TB4(2,1676,326);
    `monitor_scoreboard_upstream_connection_TB4(2,1677,327);
    `monitor_scoreboard_upstream_connection_TB4(2,1678,328);
    `monitor_scoreboard_upstream_connection_TB4(2,1679,329);
    `monitor_scoreboard_upstream_connection_TB4(2,1680,330);
    `monitor_scoreboard_upstream_connection_TB4(2,1681,331);
    `monitor_scoreboard_upstream_connection_TB4(2,1682,332);
    `monitor_scoreboard_upstream_connection_TB4(2,1683,333);
    `monitor_scoreboard_upstream_connection_TB4(2,1684,334);
    `monitor_scoreboard_upstream_connection_TB4(2,1685,335);
    `monitor_scoreboard_upstream_connection_TB4(2,1686,336);
    `monitor_scoreboard_upstream_connection_TB4(2,1687,337);
    `monitor_scoreboard_upstream_connection_TB4(2,1688,338);
    `monitor_scoreboard_upstream_connection_TB4(2,1689,339);
    `monitor_scoreboard_upstream_connection_TB4(2,1690,340);
    `monitor_scoreboard_upstream_connection_TB4(2,1691,341);
    `monitor_scoreboard_upstream_connection_TB4(2,1692,342);
    `monitor_scoreboard_upstream_connection_TB4(2,1693,343);
    `monitor_scoreboard_upstream_connection_TB4(2,1694,344);
    `monitor_scoreboard_upstream_connection_TB4(2,1695,345);
    `monitor_scoreboard_upstream_connection_TB4(2,1696,346);
    `monitor_scoreboard_upstream_connection_TB4(2,1697,347);
    `monitor_scoreboard_upstream_connection_TB4(2,1698,348);
    `monitor_scoreboard_upstream_connection_TB4(2,1699,349);
    `monitor_scoreboard_upstream_connection_TB4(2,1700,350);
    `monitor_scoreboard_upstream_connection_TB4(2,1701,351);
    `monitor_scoreboard_upstream_connection_TB4(2,1702,352);
    `monitor_scoreboard_upstream_connection_TB4(2,1703,353);
    `monitor_scoreboard_upstream_connection_TB4(2,1704,354);
    `monitor_scoreboard_upstream_connection_TB4(2,1705,355);
    `monitor_scoreboard_upstream_connection_TB4(2,1706,356);
    `monitor_scoreboard_upstream_connection_TB4(2,1707,357);
    `monitor_scoreboard_upstream_connection_TB4(2,1708,358);
    `monitor_scoreboard_upstream_connection_TB4(2,1709,359);
    `monitor_scoreboard_upstream_connection_TB4(2,1710,360);
    `monitor_scoreboard_upstream_connection_TB4(2,1711,361);
    `monitor_scoreboard_upstream_connection_TB4(2,1712,362);
    `monitor_scoreboard_upstream_connection_TB4(2,1713,363);
    `monitor_scoreboard_upstream_connection_TB4(2,1714,364);
    `monitor_scoreboard_upstream_connection_TB4(2,1715,365);
    `monitor_scoreboard_upstream_connection_TB4(2,1716,366);
    `monitor_scoreboard_upstream_connection_TB4(2,1717,367);
    `monitor_scoreboard_upstream_connection_TB4(2,1718,368);
    `monitor_scoreboard_upstream_connection_TB4(2,1719,369);
    `monitor_scoreboard_upstream_connection_TB4(2,1720,370);
    `monitor_scoreboard_upstream_connection_TB4(2,1721,371);
    `monitor_scoreboard_upstream_connection_TB4(2,1722,372);
    `monitor_scoreboard_upstream_connection_TB4(2,1723,373);
    `monitor_scoreboard_upstream_connection_TB4(2,1724,374);
    `monitor_scoreboard_upstream_connection_TB4(2,1725,375);
    `monitor_scoreboard_upstream_connection_TB4(2,1726,376);
    `monitor_scoreboard_upstream_connection_TB4(2,1727,377);
    `monitor_scoreboard_upstream_connection_TB4(2,1728,378);
    `monitor_scoreboard_upstream_connection_TB4(2,1729,379);
    `monitor_scoreboard_upstream_connection_TB4(2,1730,380);
    `monitor_scoreboard_upstream_connection_TB4(2,1731,381);
    `monitor_scoreboard_upstream_connection_TB4(2,1732,382);
    `monitor_scoreboard_upstream_connection_TB4(2,1733,383);
    `monitor_scoreboard_upstream_connection_TB4(2,1734,384);
    `monitor_scoreboard_upstream_connection_TB4(2,1735,385);
    `monitor_scoreboard_upstream_connection_TB4(2,1736,386);
    `monitor_scoreboard_upstream_connection_TB4(2,1737,387);
    `monitor_scoreboard_upstream_connection_TB4(2,1738,388);
    `monitor_scoreboard_upstream_connection_TB4(2,1739,389);
    `monitor_scoreboard_upstream_connection_TB4(2,1740,390);
    `monitor_scoreboard_upstream_connection_TB4(2,1741,391);
    `monitor_scoreboard_upstream_connection_TB4(2,1742,392);
    `monitor_scoreboard_upstream_connection_TB4(2,1743,393);
    `monitor_scoreboard_upstream_connection_TB4(2,1744,394);
    `monitor_scoreboard_upstream_connection_TB4(2,1745,395);
    `monitor_scoreboard_upstream_connection_TB4(2,1746,396);
    `monitor_scoreboard_upstream_connection_TB4(2,1747,397);
    `monitor_scoreboard_upstream_connection_TB4(2,1748,398);
    `monitor_scoreboard_upstream_connection_TB4(2,1749,399);
    `monitor_scoreboard_upstream_connection_TB4(2,1750,400);
    `monitor_scoreboard_upstream_connection_TB4(2,1751,401);
    `monitor_scoreboard_upstream_connection_TB4(2,1752,402);
    `monitor_scoreboard_upstream_connection_TB4(2,1753,403);
    `monitor_scoreboard_upstream_connection_TB4(2,1754,404);
    `monitor_scoreboard_upstream_connection_TB4(2,1755,405);
    `monitor_scoreboard_upstream_connection_TB4(2,1756,406);
    `monitor_scoreboard_upstream_connection_TB4(2,1757,407);
    `monitor_scoreboard_upstream_connection_TB4(2,1758,408);
    `monitor_scoreboard_upstream_connection_TB4(2,1759,409);
    `monitor_scoreboard_upstream_connection_TB4(2,1760,410);
    `monitor_scoreboard_upstream_connection_TB4(2,1761,411);
    `monitor_scoreboard_upstream_connection_TB4(2,1762,412);
    `monitor_scoreboard_upstream_connection_TB4(2,1763,413);
    `monitor_scoreboard_upstream_connection_TB4(2,1764,414);
    `monitor_scoreboard_upstream_connection_TB4(2,1765,415);
    `monitor_scoreboard_upstream_connection_TB4(2,1766,416);
    `monitor_scoreboard_upstream_connection_TB4(2,1767,417);
    `monitor_scoreboard_upstream_connection_TB4(2,1768,418);
    `monitor_scoreboard_upstream_connection_TB4(2,1769,419);
    `monitor_scoreboard_upstream_connection_TB4(2,1770,420);
    `monitor_scoreboard_upstream_connection_TB4(2,1771,421);
    `monitor_scoreboard_upstream_connection_TB4(2,1772,422);
    `monitor_scoreboard_upstream_connection_TB4(2,1773,423);
    `monitor_scoreboard_upstream_connection_TB4(2,1774,424);
    `monitor_scoreboard_upstream_connection_TB4(2,1775,425);
    `monitor_scoreboard_upstream_connection_TB4(2,1776,426);
    `monitor_scoreboard_upstream_connection_TB4(2,1777,427);
    `monitor_scoreboard_upstream_connection_TB4(2,1778,428);
    `monitor_scoreboard_upstream_connection_TB4(2,1779,429);
    `monitor_scoreboard_upstream_connection_TB4(2,1780,430);
    `monitor_scoreboard_upstream_connection_TB4(2,1781,431);
    `monitor_scoreboard_upstream_connection_TB4(2,1782,432);
    `monitor_scoreboard_upstream_connection_TB4(2,1783,433);
    `monitor_scoreboard_upstream_connection_TB4(2,1784,434);
    `monitor_scoreboard_upstream_connection_TB4(2,1785,435);
    `monitor_scoreboard_upstream_connection_TB4(2,1786,436);
    `monitor_scoreboard_upstream_connection_TB4(2,1787,437);
    `monitor_scoreboard_upstream_connection_TB4(2,1788,438);
    `monitor_scoreboard_upstream_connection_TB4(2,1789,439);
    `monitor_scoreboard_upstream_connection_TB4(2,1790,440);
    `monitor_scoreboard_upstream_connection_TB4(2,1791,441);
    `monitor_scoreboard_upstream_connection_TB4(2,1792,442);
    `monitor_scoreboard_upstream_connection_TB4(2,1793,443);
    `monitor_scoreboard_upstream_connection_TB4(2,1794,444);
    `monitor_scoreboard_upstream_connection_TB4(2,1795,445);
    `monitor_scoreboard_upstream_connection_TB4(2,1796,446);
    `monitor_scoreboard_upstream_connection_TB4(2,1797,447);
    `monitor_scoreboard_upstream_connection_TB4(2,1798,448);
    `monitor_scoreboard_upstream_connection_TB4(2,1799,449);
    `monitor_scoreboard_upstream_connection_TB4(3,1800,0);
    `monitor_scoreboard_upstream_connection_TB4(3,1801,1);
    `monitor_scoreboard_upstream_connection_TB4(3,1802,2);
    `monitor_scoreboard_upstream_connection_TB4(3,1803,3);
    `monitor_scoreboard_upstream_connection_TB4(3,1804,4);
    `monitor_scoreboard_upstream_connection_TB4(3,1805,5);
    `monitor_scoreboard_upstream_connection_TB4(3,1806,6);
    `monitor_scoreboard_upstream_connection_TB4(3,1807,7);
    `monitor_scoreboard_upstream_connection_TB4(3,1808,8);
    `monitor_scoreboard_upstream_connection_TB4(3,1809,9);
    `monitor_scoreboard_upstream_connection_TB4(3,1810,10);
    `monitor_scoreboard_upstream_connection_TB4(3,1811,11);
    `monitor_scoreboard_upstream_connection_TB4(3,1812,12);
    `monitor_scoreboard_upstream_connection_TB4(3,1813,13);
    `monitor_scoreboard_upstream_connection_TB4(3,1814,14);
    `monitor_scoreboard_upstream_connection_TB4(3,1815,15);
    `monitor_scoreboard_upstream_connection_TB4(3,1816,16);
    `monitor_scoreboard_upstream_connection_TB4(3,1817,17);
    `monitor_scoreboard_upstream_connection_TB4(3,1818,18);
    `monitor_scoreboard_upstream_connection_TB4(3,1819,19);
    `monitor_scoreboard_upstream_connection_TB4(3,1820,20);
    `monitor_scoreboard_upstream_connection_TB4(3,1821,21);
    `monitor_scoreboard_upstream_connection_TB4(3,1822,22);
    `monitor_scoreboard_upstream_connection_TB4(3,1823,23);
    `monitor_scoreboard_upstream_connection_TB4(3,1824,24);
    `monitor_scoreboard_upstream_connection_TB4(3,1825,25);
    `monitor_scoreboard_upstream_connection_TB4(3,1826,26);
    `monitor_scoreboard_upstream_connection_TB4(3,1827,27);
    `monitor_scoreboard_upstream_connection_TB4(3,1828,28);
    `monitor_scoreboard_upstream_connection_TB4(3,1829,29);
    `monitor_scoreboard_upstream_connection_TB4(3,1830,30);
    `monitor_scoreboard_upstream_connection_TB4(3,1831,31);
    `monitor_scoreboard_upstream_connection_TB4(3,1832,32);
    `monitor_scoreboard_upstream_connection_TB4(3,1833,33);
    `monitor_scoreboard_upstream_connection_TB4(3,1834,34);
    `monitor_scoreboard_upstream_connection_TB4(3,1835,35);
    `monitor_scoreboard_upstream_connection_TB4(3,1836,36);
    `monitor_scoreboard_upstream_connection_TB4(3,1837,37);
    `monitor_scoreboard_upstream_connection_TB4(3,1838,38);
    `monitor_scoreboard_upstream_connection_TB4(3,1839,39);
    `monitor_scoreboard_upstream_connection_TB4(3,1840,40);
    `monitor_scoreboard_upstream_connection_TB4(3,1841,41);
    `monitor_scoreboard_upstream_connection_TB4(3,1842,42);
    `monitor_scoreboard_upstream_connection_TB4(3,1843,43);
    `monitor_scoreboard_upstream_connection_TB4(3,1844,44);
    `monitor_scoreboard_upstream_connection_TB4(3,1845,45);
    `monitor_scoreboard_upstream_connection_TB4(3,1846,46);
    `monitor_scoreboard_upstream_connection_TB4(3,1847,47);
    `monitor_scoreboard_upstream_connection_TB4(3,1848,48);
    `monitor_scoreboard_upstream_connection_TB4(3,1849,49);
    `monitor_scoreboard_upstream_connection_TB4(3,1850,50);
    `monitor_scoreboard_upstream_connection_TB4(3,1851,51);
    `monitor_scoreboard_upstream_connection_TB4(3,1852,52);
    `monitor_scoreboard_upstream_connection_TB4(3,1853,53);
    `monitor_scoreboard_upstream_connection_TB4(3,1854,54);
    `monitor_scoreboard_upstream_connection_TB4(3,1855,55);
    `monitor_scoreboard_upstream_connection_TB4(3,1856,56);
    `monitor_scoreboard_upstream_connection_TB4(3,1857,57);
    `monitor_scoreboard_upstream_connection_TB4(3,1858,58);
    `monitor_scoreboard_upstream_connection_TB4(3,1859,59);
    `monitor_scoreboard_upstream_connection_TB4(3,1860,60);
    `monitor_scoreboard_upstream_connection_TB4(3,1861,61);
    `monitor_scoreboard_upstream_connection_TB4(3,1862,62);
    `monitor_scoreboard_upstream_connection_TB4(3,1863,63);
    `monitor_scoreboard_upstream_connection_TB4(3,1864,64);
    `monitor_scoreboard_upstream_connection_TB4(3,1865,65);
    `monitor_scoreboard_upstream_connection_TB4(3,1866,66);
    `monitor_scoreboard_upstream_connection_TB4(3,1867,67);
    `monitor_scoreboard_upstream_connection_TB4(3,1868,68);
    `monitor_scoreboard_upstream_connection_TB4(3,1869,69);
    `monitor_scoreboard_upstream_connection_TB4(3,1870,70);
    `monitor_scoreboard_upstream_connection_TB4(3,1871,71);
    `monitor_scoreboard_upstream_connection_TB4(3,1872,72);
    `monitor_scoreboard_upstream_connection_TB4(3,1873,73);
    `monitor_scoreboard_upstream_connection_TB4(3,1874,74);
    `monitor_scoreboard_upstream_connection_TB4(3,1875,75);
    `monitor_scoreboard_upstream_connection_TB4(3,1876,76);
    `monitor_scoreboard_upstream_connection_TB4(3,1877,77);
    `monitor_scoreboard_upstream_connection_TB4(3,1878,78);
    `monitor_scoreboard_upstream_connection_TB4(3,1879,79);
    `monitor_scoreboard_upstream_connection_TB4(3,1880,80);
    `monitor_scoreboard_upstream_connection_TB4(3,1881,81);
    `monitor_scoreboard_upstream_connection_TB4(3,1882,82);
    `monitor_scoreboard_upstream_connection_TB4(3,1883,83);
    `monitor_scoreboard_upstream_connection_TB4(3,1884,84);
    `monitor_scoreboard_upstream_connection_TB4(3,1885,85);
    `monitor_scoreboard_upstream_connection_TB4(3,1886,86);
    `monitor_scoreboard_upstream_connection_TB4(3,1887,87);
    `monitor_scoreboard_upstream_connection_TB4(3,1888,88);
    `monitor_scoreboard_upstream_connection_TB4(3,1889,89);
    `monitor_scoreboard_upstream_connection_TB4(3,1890,90);
    `monitor_scoreboard_upstream_connection_TB4(3,1891,91);
    `monitor_scoreboard_upstream_connection_TB4(3,1892,92);
    `monitor_scoreboard_upstream_connection_TB4(3,1893,93);
    `monitor_scoreboard_upstream_connection_TB4(3,1894,94);
    `monitor_scoreboard_upstream_connection_TB4(3,1895,95);
    `monitor_scoreboard_upstream_connection_TB4(3,1896,96);
    `monitor_scoreboard_upstream_connection_TB4(3,1897,97);
    `monitor_scoreboard_upstream_connection_TB4(3,1898,98);
    `monitor_scoreboard_upstream_connection_TB4(3,1899,99);
    `monitor_scoreboard_upstream_connection_TB4(3,1900,100);
    `monitor_scoreboard_upstream_connection_TB4(3,1901,101);
    `monitor_scoreboard_upstream_connection_TB4(3,1902,102);
    `monitor_scoreboard_upstream_connection_TB4(3,1903,103);
    `monitor_scoreboard_upstream_connection_TB4(3,1904,104);
    `monitor_scoreboard_upstream_connection_TB4(3,1905,105);
    `monitor_scoreboard_upstream_connection_TB4(3,1906,106);
    `monitor_scoreboard_upstream_connection_TB4(3,1907,107);
    `monitor_scoreboard_upstream_connection_TB4(3,1908,108);
    `monitor_scoreboard_upstream_connection_TB4(3,1909,109);
    `monitor_scoreboard_upstream_connection_TB4(3,1910,110);
    `monitor_scoreboard_upstream_connection_TB4(3,1911,111);
    `monitor_scoreboard_upstream_connection_TB4(3,1912,112);
    `monitor_scoreboard_upstream_connection_TB4(3,1913,113);
    `monitor_scoreboard_upstream_connection_TB4(3,1914,114);
    `monitor_scoreboard_upstream_connection_TB4(3,1915,115);
    `monitor_scoreboard_upstream_connection_TB4(3,1916,116);
    `monitor_scoreboard_upstream_connection_TB4(3,1917,117);
    `monitor_scoreboard_upstream_connection_TB4(3,1918,118);
    `monitor_scoreboard_upstream_connection_TB4(3,1919,119);
    `monitor_scoreboard_upstream_connection_TB4(3,1920,120);
    `monitor_scoreboard_upstream_connection_TB4(3,1921,121);
    `monitor_scoreboard_upstream_connection_TB4(3,1922,122);
    `monitor_scoreboard_upstream_connection_TB4(3,1923,123);
    `monitor_scoreboard_upstream_connection_TB4(3,1924,124);
    `monitor_scoreboard_upstream_connection_TB4(3,1925,125);
    `monitor_scoreboard_upstream_connection_TB4(3,1926,126);
    `monitor_scoreboard_upstream_connection_TB4(3,1927,127);
    `monitor_scoreboard_upstream_connection_TB4(3,1928,128);
    `monitor_scoreboard_upstream_connection_TB4(3,1929,129);
    `monitor_scoreboard_upstream_connection_TB4(3,1930,130);
    `monitor_scoreboard_upstream_connection_TB4(3,1931,131);
    `monitor_scoreboard_upstream_connection_TB4(3,1932,132);
    `monitor_scoreboard_upstream_connection_TB4(3,1933,133);
    `monitor_scoreboard_upstream_connection_TB4(3,1934,134);
    `monitor_scoreboard_upstream_connection_TB4(3,1935,135);
    `monitor_scoreboard_upstream_connection_TB4(3,1936,136);
    `monitor_scoreboard_upstream_connection_TB4(3,1937,137);
    `monitor_scoreboard_upstream_connection_TB4(3,1938,138);
    `monitor_scoreboard_upstream_connection_TB4(3,1939,139);
    `monitor_scoreboard_upstream_connection_TB4(3,1940,140);
    `monitor_scoreboard_upstream_connection_TB4(3,1941,141);
    `monitor_scoreboard_upstream_connection_TB4(3,1942,142);
    `monitor_scoreboard_upstream_connection_TB4(3,1943,143);
    `monitor_scoreboard_upstream_connection_TB4(3,1944,144);
    `monitor_scoreboard_upstream_connection_TB4(3,1945,145);
    `monitor_scoreboard_upstream_connection_TB4(3,1946,146);
    `monitor_scoreboard_upstream_connection_TB4(3,1947,147);
    `monitor_scoreboard_upstream_connection_TB4(3,1948,148);
    `monitor_scoreboard_upstream_connection_TB4(3,1949,149);
    `monitor_scoreboard_upstream_connection_TB4(3,1950,150);
    `monitor_scoreboard_upstream_connection_TB4(3,1951,151);
    `monitor_scoreboard_upstream_connection_TB4(3,1952,152);
    `monitor_scoreboard_upstream_connection_TB4(3,1953,153);
    `monitor_scoreboard_upstream_connection_TB4(3,1954,154);
    `monitor_scoreboard_upstream_connection_TB4(3,1955,155);
    `monitor_scoreboard_upstream_connection_TB4(3,1956,156);
    `monitor_scoreboard_upstream_connection_TB4(3,1957,157);
    `monitor_scoreboard_upstream_connection_TB4(3,1958,158);
    `monitor_scoreboard_upstream_connection_TB4(3,1959,159);
    `monitor_scoreboard_upstream_connection_TB4(3,1960,160);
    `monitor_scoreboard_upstream_connection_TB4(3,1961,161);
    `monitor_scoreboard_upstream_connection_TB4(3,1962,162);
    `monitor_scoreboard_upstream_connection_TB4(3,1963,163);
    `monitor_scoreboard_upstream_connection_TB4(3,1964,164);
    `monitor_scoreboard_upstream_connection_TB4(3,1965,165);
    `monitor_scoreboard_upstream_connection_TB4(3,1966,166);
    `monitor_scoreboard_upstream_connection_TB4(3,1967,167);
    `monitor_scoreboard_upstream_connection_TB4(3,1968,168);
    `monitor_scoreboard_upstream_connection_TB4(3,1969,169);
    `monitor_scoreboard_upstream_connection_TB4(3,1970,170);
    `monitor_scoreboard_upstream_connection_TB4(3,1971,171);
    `monitor_scoreboard_upstream_connection_TB4(3,1972,172);
    `monitor_scoreboard_upstream_connection_TB4(3,1973,173);
    `monitor_scoreboard_upstream_connection_TB4(3,1974,174);
    `monitor_scoreboard_upstream_connection_TB4(3,1975,175);
    `monitor_scoreboard_upstream_connection_TB4(3,1976,176);
    `monitor_scoreboard_upstream_connection_TB4(3,1977,177);
    `monitor_scoreboard_upstream_connection_TB4(3,1978,178);
    `monitor_scoreboard_upstream_connection_TB4(3,1979,179);
    `monitor_scoreboard_upstream_connection_TB4(3,1980,180);
    `monitor_scoreboard_upstream_connection_TB4(3,1981,181);
    `monitor_scoreboard_upstream_connection_TB4(3,1982,182);
    `monitor_scoreboard_upstream_connection_TB4(3,1983,183);
    `monitor_scoreboard_upstream_connection_TB4(3,1984,184);
    `monitor_scoreboard_upstream_connection_TB4(3,1985,185);
    `monitor_scoreboard_upstream_connection_TB4(3,1986,186);
    `monitor_scoreboard_upstream_connection_TB4(3,1987,187);
    `monitor_scoreboard_upstream_connection_TB4(3,1988,188);
    `monitor_scoreboard_upstream_connection_TB4(3,1989,189);
    `monitor_scoreboard_upstream_connection_TB4(3,1990,190);
    `monitor_scoreboard_upstream_connection_TB4(3,1991,191);
    `monitor_scoreboard_upstream_connection_TB4(3,1992,192);
    `monitor_scoreboard_upstream_connection_TB4(3,1993,193);
    `monitor_scoreboard_upstream_connection_TB4(3,1994,194);
    `monitor_scoreboard_upstream_connection_TB4(3,1995,195);
    `monitor_scoreboard_upstream_connection_TB4(3,1996,196);
    `monitor_scoreboard_upstream_connection_TB4(3,1997,197);
    `monitor_scoreboard_upstream_connection_TB4(3,1998,198);
    `monitor_scoreboard_upstream_connection_TB4(3,1999,199);
    `monitor_scoreboard_upstream_connection_TB4(3,2000,200);
    `monitor_scoreboard_upstream_connection_TB4(3,2001,201);
    `monitor_scoreboard_upstream_connection_TB4(3,2002,202);
    `monitor_scoreboard_upstream_connection_TB4(3,2003,203);
    `monitor_scoreboard_upstream_connection_TB4(3,2004,204);
    `monitor_scoreboard_upstream_connection_TB4(3,2005,205);
    `monitor_scoreboard_upstream_connection_TB4(3,2006,206);
    `monitor_scoreboard_upstream_connection_TB4(3,2007,207);
    `monitor_scoreboard_upstream_connection_TB4(3,2008,208);
    `monitor_scoreboard_upstream_connection_TB4(3,2009,209);
    `monitor_scoreboard_upstream_connection_TB4(3,2010,210);
    `monitor_scoreboard_upstream_connection_TB4(3,2011,211);
    `monitor_scoreboard_upstream_connection_TB4(3,2012,212);
    `monitor_scoreboard_upstream_connection_TB4(3,2013,213);
    `monitor_scoreboard_upstream_connection_TB4(3,2014,214);
    `monitor_scoreboard_upstream_connection_TB4(3,2015,215);
    `monitor_scoreboard_upstream_connection_TB4(3,2016,216);
    `monitor_scoreboard_upstream_connection_TB4(3,2017,217);
    `monitor_scoreboard_upstream_connection_TB4(3,2018,218);
    `monitor_scoreboard_upstream_connection_TB4(3,2019,219);
    `monitor_scoreboard_upstream_connection_TB4(3,2020,220);
    `monitor_scoreboard_upstream_connection_TB4(3,2021,221);
    `monitor_scoreboard_upstream_connection_TB4(3,2022,222);
    `monitor_scoreboard_upstream_connection_TB4(3,2023,223);
    `monitor_scoreboard_upstream_connection_TB4(3,2024,224);
    `monitor_scoreboard_upstream_connection_TB4(3,2025,225);
    `monitor_scoreboard_upstream_connection_TB4(3,2026,226);
    `monitor_scoreboard_upstream_connection_TB4(3,2027,227);
    `monitor_scoreboard_upstream_connection_TB4(3,2028,228);
    `monitor_scoreboard_upstream_connection_TB4(3,2029,229);
    `monitor_scoreboard_upstream_connection_TB4(3,2030,230);
    `monitor_scoreboard_upstream_connection_TB4(3,2031,231);
    `monitor_scoreboard_upstream_connection_TB4(3,2032,232);
    `monitor_scoreboard_upstream_connection_TB4(3,2033,233);
    `monitor_scoreboard_upstream_connection_TB4(3,2034,234);
    `monitor_scoreboard_upstream_connection_TB4(3,2035,235);
    `monitor_scoreboard_upstream_connection_TB4(3,2036,236);
    `monitor_scoreboard_upstream_connection_TB4(3,2037,237);
    `monitor_scoreboard_upstream_connection_TB4(3,2038,238);
    `monitor_scoreboard_upstream_connection_TB4(3,2039,239);
    `monitor_scoreboard_upstream_connection_TB4(3,2040,240);
    `monitor_scoreboard_upstream_connection_TB4(3,2041,241);
    `monitor_scoreboard_upstream_connection_TB4(3,2042,242);
    `monitor_scoreboard_upstream_connection_TB4(3,2043,243);
    `monitor_scoreboard_upstream_connection_TB4(3,2044,244);
    `monitor_scoreboard_upstream_connection_TB4(3,2045,245);
    `monitor_scoreboard_upstream_connection_TB4(3,2046,246);
    `monitor_scoreboard_upstream_connection_TB4(3,2047,247);
    `endif

    sequencer.master_sequencer_H =  pf_vf_mux_system_env_H.master[0].sequencer;
    sequencer.master_sequencer_D0 =  pf_vf_mux_system_env_D.master[0].sequencer;
    sequencer.master_sequencer_D1 =  pf_vf_mux_system_env_D.master[1].sequencer;
    sequencer.master_sequencer_D2 =  pf_vf_mux_system_env_D.master[2].sequencer;
    sequencer.master_sequencer_D3 =  pf_vf_mux_system_env_D.master[3].sequencer;
    sequencer.master_sequencer_D4 =  pf_vf_mux_system_env_D.master[4].sequencer;
    sequencer.master_sequencer_D5 =  pf_vf_mux_system_env_D.master[5].sequencer;
    sequencer.master_sequencer_D6 =  pf_vf_mux_system_env_D.master[6].sequencer;
    sequencer.master_sequencer_D7 =  pf_vf_mux_system_env_D.master[7].sequencer;
    sequencer.master_sequencer_D8 =  pf_vf_mux_system_env_D.master[8].sequencer;
    sequencer.master_sequencer_D9 =  pf_vf_mux_system_env_D.master[9].sequencer;
    sequencer.master_sequencer_D10 =  pf_vf_mux_system_env_D.master[10].sequencer;
    sequencer.master_sequencer_D11 =  pf_vf_mux_system_env_D.master[11].sequencer;
    sequencer.master_sequencer_D12 =  pf_vf_mux_system_env_D.master[12].sequencer;
    sequencer.master_sequencer_D13 =  pf_vf_mux_system_env_D.master[13].sequencer;
    sequencer.master_sequencer_D14 =  pf_vf_mux_system_env_D.master[14].sequencer;
    sequencer.master_sequencer_D15 =  pf_vf_mux_system_env_D.master[15].sequencer;

    `ifdef TB_CONFIG_2
    sequencer.master_sequencer_DN0 =  pf_vf_mux_system_env_DN.master[0].sequencer;
    sequencer.master_sequencer_DN1 =  pf_vf_mux_system_env_DN.master[1].sequencer;
    sequencer.master_sequencer_DN2 =  pf_vf_mux_system_env_DN.master[2].sequencer;
    sequencer.master_sequencer_DN3 =  pf_vf_mux_system_env_DN.master[3].sequencer;
    sequencer.master_sequencer_DN4 =  pf_vf_mux_system_env_DN.master[4].sequencer;
    sequencer.master_sequencer_DN5 =  pf_vf_mux_system_env_DN.master[5].sequencer;
    sequencer.master_sequencer_DN6 =  pf_vf_mux_system_env_DN.master[6].sequencer;
    sequencer.master_sequencer_DN7 =  pf_vf_mux_system_env_DN.master[7].sequencer;
    `elsif TB_CONFIG_3
    sequencer.master_sequencer_DN0 =  pf_vf_mux_system_env_DN.master[0].sequencer;
    sequencer.master_sequencer_DN1 =  pf_vf_mux_system_env_DN.master[1].sequencer;
    sequencer.master_sequencer_DN2 =  pf_vf_mux_system_env_DN.master[2].sequencer;
    sequencer.master_sequencer_DN3 =  pf_vf_mux_system_env_DN.master[3].sequencer;
    sequencer.master_sequencer_DN4 =  pf_vf_mux_system_env_DN.master[4].sequencer;
    sequencer.master_sequencer_DN5 =  pf_vf_mux_system_env_DN.master[5].sequencer;
    sequencer.master_sequencer_DN6 =  pf_vf_mux_system_env_DN.master[6].sequencer;
    sequencer.master_sequencer_DN7 =  pf_vf_mux_system_env_DN.master[7].sequencer;
    sequencer.master_sequencer_DN8 =  pf_vf_mux_system_env_DN.master[8].sequencer;
    sequencer.master_sequencer_DN9 =  pf_vf_mux_system_env_DN.master[9].sequencer;
    sequencer.master_sequencer_DN10 =  pf_vf_mux_system_env_DN.master[10].sequencer;
    sequencer.master_sequencer_DN11 =  pf_vf_mux_system_env_DN.master[11].sequencer;
    sequencer.master_sequencer_DN12 =  pf_vf_mux_system_env_DN.master[12].sequencer;
    sequencer.master_sequencer_DN13 =  pf_vf_mux_system_env_DN.master[13].sequencer;
    sequencer.master_sequencer_DN14 =  pf_vf_mux_system_env_DN.master[14].sequencer;
    sequencer.master_sequencer_DN15 =  pf_vf_mux_system_env_DN.master[15].sequencer;
    `elsif TB_CONFIG_4
    sequencer.master_sequencer_D16 =  pf_vf_mux_system_env_D.master[16].sequencer;
    sequencer.master_sequencer_D17 =  pf_vf_mux_system_env_D.master[17].sequencer;
    sequencer.master_sequencer_D18 =  pf_vf_mux_system_env_D.master[18].sequencer;
    sequencer.master_sequencer_D19 =  pf_vf_mux_system_env_D.master[19].sequencer;
    sequencer.master_sequencer_D20 =  pf_vf_mux_system_env_D.master[20].sequencer;
    sequencer.master_sequencer_D21 =  pf_vf_mux_system_env_D.master[21].sequencer;
    sequencer.master_sequencer_D22 =  pf_vf_mux_system_env_D.master[22].sequencer;
    sequencer.master_sequencer_D23 =  pf_vf_mux_system_env_D.master[23].sequencer;
    sequencer.master_sequencer_D24 =  pf_vf_mux_system_env_D.master[24].sequencer;
    sequencer.master_sequencer_D25 =  pf_vf_mux_system_env_D.master[25].sequencer;
    sequencer.master_sequencer_D26 =  pf_vf_mux_system_env_D.master[26].sequencer;
    sequencer.master_sequencer_D27 =  pf_vf_mux_system_env_D.master[27].sequencer;
    sequencer.master_sequencer_D28 =  pf_vf_mux_system_env_D.master[28].sequencer;
    sequencer.master_sequencer_D29 =  pf_vf_mux_system_env_D.master[29].sequencer;
    sequencer.master_sequencer_D30 =  pf_vf_mux_system_env_D.master[30].sequencer;
    sequencer.master_sequencer_D31 =  pf_vf_mux_system_env_D.master[31].sequencer;
    sequencer.master_sequencer_D32 =  pf_vf_mux_system_env_D.master[32].sequencer;
    sequencer.master_sequencer_D33 =  pf_vf_mux_system_env_D.master[33].sequencer;
    sequencer.master_sequencer_D34 =  pf_vf_mux_system_env_D.master[34].sequencer;
    sequencer.master_sequencer_D35 =  pf_vf_mux_system_env_D.master[35].sequencer;
    sequencer.master_sequencer_D36 =  pf_vf_mux_system_env_D.master[36].sequencer;
    sequencer.master_sequencer_D37 =  pf_vf_mux_system_env_D.master[37].sequencer;
    sequencer.master_sequencer_D38 =  pf_vf_mux_system_env_D.master[38].sequencer;
    sequencer.master_sequencer_D39 =  pf_vf_mux_system_env_D.master[39].sequencer;
    sequencer.master_sequencer_D40 =  pf_vf_mux_system_env_D.master[40].sequencer;
    sequencer.master_sequencer_D41 =  pf_vf_mux_system_env_D.master[41].sequencer;
    sequencer.master_sequencer_D42 =  pf_vf_mux_system_env_D.master[42].sequencer;
    sequencer.master_sequencer_D43 =  pf_vf_mux_system_env_D.master[43].sequencer;
    sequencer.master_sequencer_D44 =  pf_vf_mux_system_env_D.master[44].sequencer;
    sequencer.master_sequencer_D45 =  pf_vf_mux_system_env_D.master[45].sequencer;
    sequencer.master_sequencer_D46 =  pf_vf_mux_system_env_D.master[46].sequencer;
    sequencer.master_sequencer_D47 =  pf_vf_mux_system_env_D.master[47].sequencer;
    sequencer.master_sequencer_D48 =  pf_vf_mux_system_env_D.master[48].sequencer;
    sequencer.master_sequencer_D49 =  pf_vf_mux_system_env_D.master[49].sequencer;
    sequencer.master_sequencer_D50 =  pf_vf_mux_system_env_D.master[50].sequencer;
    sequencer.master_sequencer_D51 =  pf_vf_mux_system_env_D.master[51].sequencer;
    sequencer.master_sequencer_D52 =  pf_vf_mux_system_env_D.master[52].sequencer;
    sequencer.master_sequencer_D53 =  pf_vf_mux_system_env_D.master[53].sequencer;
    sequencer.master_sequencer_D54 =  pf_vf_mux_system_env_D.master[54].sequencer;
    sequencer.master_sequencer_D55 =  pf_vf_mux_system_env_D.master[55].sequencer;
    sequencer.master_sequencer_D56 =  pf_vf_mux_system_env_D.master[56].sequencer;
    sequencer.master_sequencer_D57 =  pf_vf_mux_system_env_D.master[57].sequencer;
    sequencer.master_sequencer_D58 =  pf_vf_mux_system_env_D.master[58].sequencer;
    sequencer.master_sequencer_D59 =  pf_vf_mux_system_env_D.master[59].sequencer;
    sequencer.master_sequencer_D60 =  pf_vf_mux_system_env_D.master[60].sequencer;
    sequencer.master_sequencer_D61 =  pf_vf_mux_system_env_D.master[61].sequencer;
    sequencer.master_sequencer_D62 =  pf_vf_mux_system_env_D.master[62].sequencer;
    sequencer.master_sequencer_D63 =  pf_vf_mux_system_env_D.master[63].sequencer;
    sequencer.master_sequencer_D64 =  pf_vf_mux_system_env_D.master[64].sequencer;
    sequencer.master_sequencer_D65 =  pf_vf_mux_system_env_D.master[65].sequencer;
    sequencer.master_sequencer_D66 =  pf_vf_mux_system_env_D.master[66].sequencer;
    sequencer.master_sequencer_D67 =  pf_vf_mux_system_env_D.master[67].sequencer;
    sequencer.master_sequencer_D68 =  pf_vf_mux_system_env_D.master[68].sequencer;
    sequencer.master_sequencer_D69 =  pf_vf_mux_system_env_D.master[69].sequencer;
    sequencer.master_sequencer_D70 =  pf_vf_mux_system_env_D.master[70].sequencer;
    sequencer.master_sequencer_D71 =  pf_vf_mux_system_env_D.master[71].sequencer;
    sequencer.master_sequencer_D72 =  pf_vf_mux_system_env_D.master[72].sequencer;
    sequencer.master_sequencer_D73 =  pf_vf_mux_system_env_D.master[73].sequencer;
    sequencer.master_sequencer_D74 =  pf_vf_mux_system_env_D.master[74].sequencer;
    sequencer.master_sequencer_D75 =  pf_vf_mux_system_env_D.master[75].sequencer;
    sequencer.master_sequencer_D76 =  pf_vf_mux_system_env_D.master[76].sequencer;
    sequencer.master_sequencer_D77 =  pf_vf_mux_system_env_D.master[77].sequencer;
    sequencer.master_sequencer_D78 =  pf_vf_mux_system_env_D.master[78].sequencer;
    sequencer.master_sequencer_D79 =  pf_vf_mux_system_env_D.master[79].sequencer;
    sequencer.master_sequencer_D80 =  pf_vf_mux_system_env_D.master[80].sequencer;
    sequencer.master_sequencer_D81 =  pf_vf_mux_system_env_D.master[81].sequencer;
    sequencer.master_sequencer_D82 =  pf_vf_mux_system_env_D.master[82].sequencer;
    sequencer.master_sequencer_D83 =  pf_vf_mux_system_env_D.master[83].sequencer;
    sequencer.master_sequencer_D84 =  pf_vf_mux_system_env_D.master[84].sequencer;
    sequencer.master_sequencer_D85 =  pf_vf_mux_system_env_D.master[85].sequencer;
    sequencer.master_sequencer_D86 =  pf_vf_mux_system_env_D.master[86].sequencer;
    sequencer.master_sequencer_D87 =  pf_vf_mux_system_env_D.master[87].sequencer;
    sequencer.master_sequencer_D88 =  pf_vf_mux_system_env_D.master[88].sequencer;
    sequencer.master_sequencer_D89 =  pf_vf_mux_system_env_D.master[89].sequencer;
    sequencer.master_sequencer_D90 =  pf_vf_mux_system_env_D.master[90].sequencer;
    sequencer.master_sequencer_D91 =  pf_vf_mux_system_env_D.master[91].sequencer;
    sequencer.master_sequencer_D92 =  pf_vf_mux_system_env_D.master[92].sequencer;
    sequencer.master_sequencer_D93 =  pf_vf_mux_system_env_D.master[93].sequencer;
    sequencer.master_sequencer_D94 =  pf_vf_mux_system_env_D.master[94].sequencer;
    sequencer.master_sequencer_D95 =  pf_vf_mux_system_env_D.master[95].sequencer;
    sequencer.master_sequencer_D96 =  pf_vf_mux_system_env_D.master[96].sequencer;
    sequencer.master_sequencer_D97 =  pf_vf_mux_system_env_D.master[97].sequencer;
    sequencer.master_sequencer_D98 =  pf_vf_mux_system_env_D.master[98].sequencer;
    sequencer.master_sequencer_D99 =  pf_vf_mux_system_env_D.master[99].sequencer;
    sequencer.master_sequencer_D100 =  pf_vf_mux_system_env_D.master[100].sequencer;
    sequencer.master_sequencer_D101 =  pf_vf_mux_system_env_D.master[101].sequencer;
    sequencer.master_sequencer_D102 =  pf_vf_mux_system_env_D.master[102].sequencer;
    sequencer.master_sequencer_D103 =  pf_vf_mux_system_env_D.master[103].sequencer;
    sequencer.master_sequencer_D104 =  pf_vf_mux_system_env_D.master[104].sequencer;
    sequencer.master_sequencer_D105 =  pf_vf_mux_system_env_D.master[105].sequencer;
    sequencer.master_sequencer_D106 =  pf_vf_mux_system_env_D.master[106].sequencer;
    sequencer.master_sequencer_D107 =  pf_vf_mux_system_env_D.master[107].sequencer;
    sequencer.master_sequencer_D108 =  pf_vf_mux_system_env_D.master[108].sequencer;
    sequencer.master_sequencer_D109 =  pf_vf_mux_system_env_D.master[109].sequencer;
    sequencer.master_sequencer_D110 =  pf_vf_mux_system_env_D.master[110].sequencer;
    sequencer.master_sequencer_D111 =  pf_vf_mux_system_env_D.master[111].sequencer;
    sequencer.master_sequencer_D112 =  pf_vf_mux_system_env_D.master[112].sequencer;
    sequencer.master_sequencer_D113 =  pf_vf_mux_system_env_D.master[113].sequencer;
    sequencer.master_sequencer_D114 =  pf_vf_mux_system_env_D.master[114].sequencer;
    sequencer.master_sequencer_D115 =  pf_vf_mux_system_env_D.master[115].sequencer;
    sequencer.master_sequencer_D116 =  pf_vf_mux_system_env_D.master[116].sequencer;
    sequencer.master_sequencer_D117 =  pf_vf_mux_system_env_D.master[117].sequencer;
    sequencer.master_sequencer_D118 =  pf_vf_mux_system_env_D.master[118].sequencer;
    sequencer.master_sequencer_D119 =  pf_vf_mux_system_env_D.master[119].sequencer;
    sequencer.master_sequencer_D120 =  pf_vf_mux_system_env_D.master[120].sequencer;
    sequencer.master_sequencer_D121 =  pf_vf_mux_system_env_D.master[121].sequencer;
    sequencer.master_sequencer_D122 =  pf_vf_mux_system_env_D.master[122].sequencer;
    sequencer.master_sequencer_D123 =  pf_vf_mux_system_env_D.master[123].sequencer;
    sequencer.master_sequencer_D124 =  pf_vf_mux_system_env_D.master[124].sequencer;
    sequencer.master_sequencer_D125 =  pf_vf_mux_system_env_D.master[125].sequencer;
    sequencer.master_sequencer_D126 =  pf_vf_mux_system_env_D.master[126].sequencer;
    sequencer.master_sequencer_D127 =  pf_vf_mux_system_env_D.master[127].sequencer;
    sequencer.master_sequencer_D128 =  pf_vf_mux_system_env_D.master[128].sequencer;
    sequencer.master_sequencer_D129 =  pf_vf_mux_system_env_D.master[129].sequencer;
    sequencer.master_sequencer_D130 =  pf_vf_mux_system_env_D.master[130].sequencer;
    sequencer.master_sequencer_D131 =  pf_vf_mux_system_env_D.master[131].sequencer;
    sequencer.master_sequencer_D132 =  pf_vf_mux_system_env_D.master[132].sequencer;
    sequencer.master_sequencer_D133 =  pf_vf_mux_system_env_D.master[133].sequencer;
    sequencer.master_sequencer_D134 =  pf_vf_mux_system_env_D.master[134].sequencer;
    sequencer.master_sequencer_D135 =  pf_vf_mux_system_env_D.master[135].sequencer;
    sequencer.master_sequencer_D136 =  pf_vf_mux_system_env_D.master[136].sequencer;
    sequencer.master_sequencer_D137 =  pf_vf_mux_system_env_D.master[137].sequencer;
    sequencer.master_sequencer_D138 =  pf_vf_mux_system_env_D.master[138].sequencer;
    sequencer.master_sequencer_D139 =  pf_vf_mux_system_env_D.master[139].sequencer;
    sequencer.master_sequencer_D140 =  pf_vf_mux_system_env_D.master[140].sequencer;
    sequencer.master_sequencer_D141 =  pf_vf_mux_system_env_D.master[141].sequencer;
    sequencer.master_sequencer_D142 =  pf_vf_mux_system_env_D.master[142].sequencer;
    sequencer.master_sequencer_D143 =  pf_vf_mux_system_env_D.master[143].sequencer;
    sequencer.master_sequencer_D144 =  pf_vf_mux_system_env_D.master[144].sequencer;
    sequencer.master_sequencer_D145 =  pf_vf_mux_system_env_D.master[145].sequencer;
    sequencer.master_sequencer_D146 =  pf_vf_mux_system_env_D.master[146].sequencer;
    sequencer.master_sequencer_D147 =  pf_vf_mux_system_env_D.master[147].sequencer;
    sequencer.master_sequencer_D148 =  pf_vf_mux_system_env_D.master[148].sequencer;
    sequencer.master_sequencer_D149 =  pf_vf_mux_system_env_D.master[149].sequencer;
    sequencer.master_sequencer_D150 =  pf_vf_mux_system_env_D.master[150].sequencer;
    sequencer.master_sequencer_D151 =  pf_vf_mux_system_env_D.master[151].sequencer;
    sequencer.master_sequencer_D152 =  pf_vf_mux_system_env_D.master[152].sequencer;
    sequencer.master_sequencer_D153 =  pf_vf_mux_system_env_D.master[153].sequencer;
    sequencer.master_sequencer_D154 =  pf_vf_mux_system_env_D.master[154].sequencer;
    sequencer.master_sequencer_D155 =  pf_vf_mux_system_env_D.master[155].sequencer;
    sequencer.master_sequencer_D156 =  pf_vf_mux_system_env_D.master[156].sequencer;
    sequencer.master_sequencer_D157 =  pf_vf_mux_system_env_D.master[157].sequencer;
    sequencer.master_sequencer_D158 =  pf_vf_mux_system_env_D.master[158].sequencer;
    sequencer.master_sequencer_D159 =  pf_vf_mux_system_env_D.master[159].sequencer;
    sequencer.master_sequencer_D160 =  pf_vf_mux_system_env_D.master[160].sequencer;
    sequencer.master_sequencer_D161 =  pf_vf_mux_system_env_D.master[161].sequencer;
    sequencer.master_sequencer_D162 =  pf_vf_mux_system_env_D.master[162].sequencer;
    sequencer.master_sequencer_D163 =  pf_vf_mux_system_env_D.master[163].sequencer;
    sequencer.master_sequencer_D164 =  pf_vf_mux_system_env_D.master[164].sequencer;
    sequencer.master_sequencer_D165 =  pf_vf_mux_system_env_D.master[165].sequencer;
    sequencer.master_sequencer_D166 =  pf_vf_mux_system_env_D.master[166].sequencer;
    sequencer.master_sequencer_D167 =  pf_vf_mux_system_env_D.master[167].sequencer;
    sequencer.master_sequencer_D168 =  pf_vf_mux_system_env_D.master[168].sequencer;
    sequencer.master_sequencer_D169 =  pf_vf_mux_system_env_D.master[169].sequencer;
    sequencer.master_sequencer_D170 =  pf_vf_mux_system_env_D.master[170].sequencer;
    sequencer.master_sequencer_D171 =  pf_vf_mux_system_env_D.master[171].sequencer;
    sequencer.master_sequencer_D172 =  pf_vf_mux_system_env_D.master[172].sequencer;
    sequencer.master_sequencer_D173 =  pf_vf_mux_system_env_D.master[173].sequencer;
    sequencer.master_sequencer_D174 =  pf_vf_mux_system_env_D.master[174].sequencer;
    sequencer.master_sequencer_D175 =  pf_vf_mux_system_env_D.master[175].sequencer;
    sequencer.master_sequencer_D176 =  pf_vf_mux_system_env_D.master[176].sequencer;
    sequencer.master_sequencer_D177 =  pf_vf_mux_system_env_D.master[177].sequencer;
    sequencer.master_sequencer_D178 =  pf_vf_mux_system_env_D.master[178].sequencer;
    sequencer.master_sequencer_D179 =  pf_vf_mux_system_env_D.master[179].sequencer;
    sequencer.master_sequencer_D180 =  pf_vf_mux_system_env_D.master[180].sequencer;
    sequencer.master_sequencer_D181 =  pf_vf_mux_system_env_D.master[181].sequencer;
    sequencer.master_sequencer_D182 =  pf_vf_mux_system_env_D.master[182].sequencer;
    sequencer.master_sequencer_D183 =  pf_vf_mux_system_env_D.master[183].sequencer;
    sequencer.master_sequencer_D184 =  pf_vf_mux_system_env_D.master[184].sequencer;
    sequencer.master_sequencer_D185 =  pf_vf_mux_system_env_D.master[185].sequencer;
    sequencer.master_sequencer_D186 =  pf_vf_mux_system_env_D.master[186].sequencer;
    sequencer.master_sequencer_D187 =  pf_vf_mux_system_env_D.master[187].sequencer;
    sequencer.master_sequencer_D188 =  pf_vf_mux_system_env_D.master[188].sequencer;
    sequencer.master_sequencer_D189 =  pf_vf_mux_system_env_D.master[189].sequencer;
    sequencer.master_sequencer_D190 =  pf_vf_mux_system_env_D.master[190].sequencer;
    sequencer.master_sequencer_D191 =  pf_vf_mux_system_env_D.master[191].sequencer;
    sequencer.master_sequencer_D192 =  pf_vf_mux_system_env_D.master[192].sequencer;
    sequencer.master_sequencer_D193 =  pf_vf_mux_system_env_D.master[193].sequencer;
    sequencer.master_sequencer_D194 =  pf_vf_mux_system_env_D.master[194].sequencer;
    sequencer.master_sequencer_D195 =  pf_vf_mux_system_env_D.master[195].sequencer;
    sequencer.master_sequencer_D196 =  pf_vf_mux_system_env_D.master[196].sequencer;
    sequencer.master_sequencer_D197 =  pf_vf_mux_system_env_D.master[197].sequencer;
    sequencer.master_sequencer_D198 =  pf_vf_mux_system_env_D.master[198].sequencer;
    sequencer.master_sequencer_D199 =  pf_vf_mux_system_env_D.master[199].sequencer;
    sequencer.master_sequencer_D200 =  pf_vf_mux_system_env_D.master[200].sequencer;
    sequencer.master_sequencer_D201 =  pf_vf_mux_system_env_D.master[201].sequencer;
    sequencer.master_sequencer_D202 =  pf_vf_mux_system_env_D.master[202].sequencer;
    sequencer.master_sequencer_D203 =  pf_vf_mux_system_env_D.master[203].sequencer;
    sequencer.master_sequencer_D204 =  pf_vf_mux_system_env_D.master[204].sequencer;
    sequencer.master_sequencer_D205 =  pf_vf_mux_system_env_D.master[205].sequencer;
    sequencer.master_sequencer_D206 =  pf_vf_mux_system_env_D.master[206].sequencer;
    sequencer.master_sequencer_D207 =  pf_vf_mux_system_env_D.master[207].sequencer;
    sequencer.master_sequencer_D208 =  pf_vf_mux_system_env_D.master[208].sequencer;
    sequencer.master_sequencer_D209 =  pf_vf_mux_system_env_D.master[209].sequencer;
    sequencer.master_sequencer_D210 =  pf_vf_mux_system_env_D.master[210].sequencer;
    sequencer.master_sequencer_D211 =  pf_vf_mux_system_env_D.master[211].sequencer;
    sequencer.master_sequencer_D212 =  pf_vf_mux_system_env_D.master[212].sequencer;
    sequencer.master_sequencer_D213 =  pf_vf_mux_system_env_D.master[213].sequencer;
    sequencer.master_sequencer_D214 =  pf_vf_mux_system_env_D.master[214].sequencer;
    sequencer.master_sequencer_D215 =  pf_vf_mux_system_env_D.master[215].sequencer;
    sequencer.master_sequencer_D216 =  pf_vf_mux_system_env_D.master[216].sequencer;
    sequencer.master_sequencer_D217 =  pf_vf_mux_system_env_D.master[217].sequencer;
    sequencer.master_sequencer_D218 =  pf_vf_mux_system_env_D.master[218].sequencer;
    sequencer.master_sequencer_D219 =  pf_vf_mux_system_env_D.master[219].sequencer;
    sequencer.master_sequencer_D220 =  pf_vf_mux_system_env_D.master[220].sequencer;
    sequencer.master_sequencer_D221 =  pf_vf_mux_system_env_D.master[221].sequencer;
    sequencer.master_sequencer_D222 =  pf_vf_mux_system_env_D.master[222].sequencer;
    sequencer.master_sequencer_D223 =  pf_vf_mux_system_env_D.master[223].sequencer;
    sequencer.master_sequencer_D224 =  pf_vf_mux_system_env_D.master[224].sequencer;
    sequencer.master_sequencer_D225 =  pf_vf_mux_system_env_D.master[225].sequencer;
    sequencer.master_sequencer_D226 =  pf_vf_mux_system_env_D.master[226].sequencer;
    sequencer.master_sequencer_D227 =  pf_vf_mux_system_env_D.master[227].sequencer;
    sequencer.master_sequencer_D228 =  pf_vf_mux_system_env_D.master[228].sequencer;
    sequencer.master_sequencer_D229 =  pf_vf_mux_system_env_D.master[229].sequencer;
    sequencer.master_sequencer_D230 =  pf_vf_mux_system_env_D.master[230].sequencer;
    sequencer.master_sequencer_D231 =  pf_vf_mux_system_env_D.master[231].sequencer;
    sequencer.master_sequencer_D232 =  pf_vf_mux_system_env_D.master[232].sequencer;
    sequencer.master_sequencer_D233 =  pf_vf_mux_system_env_D.master[233].sequencer;
    sequencer.master_sequencer_D234 =  pf_vf_mux_system_env_D.master[234].sequencer;
    sequencer.master_sequencer_D235 =  pf_vf_mux_system_env_D.master[235].sequencer;
    sequencer.master_sequencer_D236 =  pf_vf_mux_system_env_D.master[236].sequencer;
    sequencer.master_sequencer_D237 =  pf_vf_mux_system_env_D.master[237].sequencer;
    sequencer.master_sequencer_D238 =  pf_vf_mux_system_env_D.master[238].sequencer;
    sequencer.master_sequencer_D239 =  pf_vf_mux_system_env_D.master[239].sequencer;
    sequencer.master_sequencer_D240 =  pf_vf_mux_system_env_D.master[240].sequencer;
    sequencer.master_sequencer_D241 =  pf_vf_mux_system_env_D.master[241].sequencer;
    sequencer.master_sequencer_D242 =  pf_vf_mux_system_env_D.master[242].sequencer;
    sequencer.master_sequencer_D243 =  pf_vf_mux_system_env_D.master[243].sequencer;
    sequencer.master_sequencer_D244 =  pf_vf_mux_system_env_D.master[244].sequencer;
    sequencer.master_sequencer_D245 =  pf_vf_mux_system_env_D.master[245].sequencer;
    sequencer.master_sequencer_D246 =  pf_vf_mux_system_env_D.master[246].sequencer;
    sequencer.master_sequencer_D247 =  pf_vf_mux_system_env_D.master[247].sequencer;
    sequencer.master_sequencer_D248 =  pf_vf_mux_system_env_D.master[248].sequencer;
    sequencer.master_sequencer_D249 =  pf_vf_mux_system_env_D.master[249].sequencer;
    sequencer.master_sequencer_D250 =  pf_vf_mux_system_env_D.master[250].sequencer;
    sequencer.master_sequencer_D251 =  pf_vf_mux_system_env_D.master[251].sequencer;
    sequencer.master_sequencer_D252 =  pf_vf_mux_system_env_D.master[252].sequencer;
    sequencer.master_sequencer_D253 =  pf_vf_mux_system_env_D.master[253].sequencer;
    sequencer.master_sequencer_D254 =  pf_vf_mux_system_env_D.master[254].sequencer;
    sequencer.master_sequencer_D255 =  pf_vf_mux_system_env_D.master[255].sequencer;
    sequencer.master_sequencer_D256 =  pf_vf_mux_system_env_D.master[256].sequencer;
    sequencer.master_sequencer_D257 =  pf_vf_mux_system_env_D.master[257].sequencer;
    sequencer.master_sequencer_D258 =  pf_vf_mux_system_env_D.master[258].sequencer;
    sequencer.master_sequencer_D259 =  pf_vf_mux_system_env_D.master[259].sequencer;
    sequencer.master_sequencer_D260 =  pf_vf_mux_system_env_D.master[260].sequencer;
    sequencer.master_sequencer_D261 =  pf_vf_mux_system_env_D.master[261].sequencer;
    sequencer.master_sequencer_D262 =  pf_vf_mux_system_env_D.master[262].sequencer;
    sequencer.master_sequencer_D263 =  pf_vf_mux_system_env_D.master[263].sequencer;
    sequencer.master_sequencer_D264 =  pf_vf_mux_system_env_D.master[264].sequencer;
    sequencer.master_sequencer_D265 =  pf_vf_mux_system_env_D.master[265].sequencer;
    sequencer.master_sequencer_D266 =  pf_vf_mux_system_env_D.master[266].sequencer;
    sequencer.master_sequencer_D267 =  pf_vf_mux_system_env_D.master[267].sequencer;
    sequencer.master_sequencer_D268 =  pf_vf_mux_system_env_D.master[268].sequencer;
    sequencer.master_sequencer_D269 =  pf_vf_mux_system_env_D.master[269].sequencer;
    sequencer.master_sequencer_D270 =  pf_vf_mux_system_env_D.master[270].sequencer;
    sequencer.master_sequencer_D271 =  pf_vf_mux_system_env_D.master[271].sequencer;
    sequencer.master_sequencer_D272 =  pf_vf_mux_system_env_D.master[272].sequencer;
    sequencer.master_sequencer_D273 =  pf_vf_mux_system_env_D.master[273].sequencer;
    sequencer.master_sequencer_D274 =  pf_vf_mux_system_env_D.master[274].sequencer;
    sequencer.master_sequencer_D275 =  pf_vf_mux_system_env_D.master[275].sequencer;
    sequencer.master_sequencer_D276 =  pf_vf_mux_system_env_D.master[276].sequencer;
    sequencer.master_sequencer_D277 =  pf_vf_mux_system_env_D.master[277].sequencer;
    sequencer.master_sequencer_D278 =  pf_vf_mux_system_env_D.master[278].sequencer;
    sequencer.master_sequencer_D279 =  pf_vf_mux_system_env_D.master[279].sequencer;
    sequencer.master_sequencer_D280 =  pf_vf_mux_system_env_D.master[280].sequencer;
    sequencer.master_sequencer_D281 =  pf_vf_mux_system_env_D.master[281].sequencer;
    sequencer.master_sequencer_D282 =  pf_vf_mux_system_env_D.master[282].sequencer;
    sequencer.master_sequencer_D283 =  pf_vf_mux_system_env_D.master[283].sequencer;
    sequencer.master_sequencer_D284 =  pf_vf_mux_system_env_D.master[284].sequencer;
    sequencer.master_sequencer_D285 =  pf_vf_mux_system_env_D.master[285].sequencer;
    sequencer.master_sequencer_D286 =  pf_vf_mux_system_env_D.master[286].sequencer;
    sequencer.master_sequencer_D287 =  pf_vf_mux_system_env_D.master[287].sequencer;
    sequencer.master_sequencer_D288 =  pf_vf_mux_system_env_D.master[288].sequencer;
    sequencer.master_sequencer_D289 =  pf_vf_mux_system_env_D.master[289].sequencer;
    sequencer.master_sequencer_D290 =  pf_vf_mux_system_env_D.master[290].sequencer;
    sequencer.master_sequencer_D291 =  pf_vf_mux_system_env_D.master[291].sequencer;
    sequencer.master_sequencer_D292 =  pf_vf_mux_system_env_D.master[292].sequencer;
    sequencer.master_sequencer_D293 =  pf_vf_mux_system_env_D.master[293].sequencer;
    sequencer.master_sequencer_D294 =  pf_vf_mux_system_env_D.master[294].sequencer;
    sequencer.master_sequencer_D295 =  pf_vf_mux_system_env_D.master[295].sequencer;
    sequencer.master_sequencer_D296 =  pf_vf_mux_system_env_D.master[296].sequencer;
    sequencer.master_sequencer_D297 =  pf_vf_mux_system_env_D.master[297].sequencer;
    sequencer.master_sequencer_D298 =  pf_vf_mux_system_env_D.master[298].sequencer;
    sequencer.master_sequencer_D299 =  pf_vf_mux_system_env_D.master[299].sequencer;
    sequencer.master_sequencer_D300 =  pf_vf_mux_system_env_D.master[300].sequencer;
    sequencer.master_sequencer_D301 =  pf_vf_mux_system_env_D.master[301].sequencer;
    sequencer.master_sequencer_D302 =  pf_vf_mux_system_env_D.master[302].sequencer;
    sequencer.master_sequencer_D303 =  pf_vf_mux_system_env_D.master[303].sequencer;
    sequencer.master_sequencer_D304 =  pf_vf_mux_system_env_D.master[304].sequencer;
    sequencer.master_sequencer_D305 =  pf_vf_mux_system_env_D.master[305].sequencer;
    sequencer.master_sequencer_D306 =  pf_vf_mux_system_env_D.master[306].sequencer;
    sequencer.master_sequencer_D307 =  pf_vf_mux_system_env_D.master[307].sequencer;
    sequencer.master_sequencer_D308 =  pf_vf_mux_system_env_D.master[308].sequencer;
    sequencer.master_sequencer_D309 =  pf_vf_mux_system_env_D.master[309].sequencer;
    sequencer.master_sequencer_D310 =  pf_vf_mux_system_env_D.master[310].sequencer;
    sequencer.master_sequencer_D311 =  pf_vf_mux_system_env_D.master[311].sequencer;
    sequencer.master_sequencer_D312 =  pf_vf_mux_system_env_D.master[312].sequencer;
    sequencer.master_sequencer_D313 =  pf_vf_mux_system_env_D.master[313].sequencer;
    sequencer.master_sequencer_D314 =  pf_vf_mux_system_env_D.master[314].sequencer;
    sequencer.master_sequencer_D315 =  pf_vf_mux_system_env_D.master[315].sequencer;
    sequencer.master_sequencer_D316 =  pf_vf_mux_system_env_D.master[316].sequencer;
    sequencer.master_sequencer_D317 =  pf_vf_mux_system_env_D.master[317].sequencer;
    sequencer.master_sequencer_D318 =  pf_vf_mux_system_env_D.master[318].sequencer;
    sequencer.master_sequencer_D319 =  pf_vf_mux_system_env_D.master[319].sequencer;
    sequencer.master_sequencer_D320 =  pf_vf_mux_system_env_D.master[320].sequencer;
    sequencer.master_sequencer_D321 =  pf_vf_mux_system_env_D.master[321].sequencer;
    sequencer.master_sequencer_D322 =  pf_vf_mux_system_env_D.master[322].sequencer;
    sequencer.master_sequencer_D323 =  pf_vf_mux_system_env_D.master[323].sequencer;
    sequencer.master_sequencer_D324 =  pf_vf_mux_system_env_D.master[324].sequencer;
    sequencer.master_sequencer_D325 =  pf_vf_mux_system_env_D.master[325].sequencer;
    sequencer.master_sequencer_D326 =  pf_vf_mux_system_env_D.master[326].sequencer;
    sequencer.master_sequencer_D327 =  pf_vf_mux_system_env_D.master[327].sequencer;
    sequencer.master_sequencer_D328 =  pf_vf_mux_system_env_D.master[328].sequencer;
    sequencer.master_sequencer_D329 =  pf_vf_mux_system_env_D.master[329].sequencer;
    sequencer.master_sequencer_D330 =  pf_vf_mux_system_env_D.master[330].sequencer;
    sequencer.master_sequencer_D331 =  pf_vf_mux_system_env_D.master[331].sequencer;
    sequencer.master_sequencer_D332 =  pf_vf_mux_system_env_D.master[332].sequencer;
    sequencer.master_sequencer_D333 =  pf_vf_mux_system_env_D.master[333].sequencer;
    sequencer.master_sequencer_D334 =  pf_vf_mux_system_env_D.master[334].sequencer;
    sequencer.master_sequencer_D335 =  pf_vf_mux_system_env_D.master[335].sequencer;
    sequencer.master_sequencer_D336 =  pf_vf_mux_system_env_D.master[336].sequencer;
    sequencer.master_sequencer_D337 =  pf_vf_mux_system_env_D.master[337].sequencer;
    sequencer.master_sequencer_D338 =  pf_vf_mux_system_env_D.master[338].sequencer;
    sequencer.master_sequencer_D339 =  pf_vf_mux_system_env_D.master[339].sequencer;
    sequencer.master_sequencer_D340 =  pf_vf_mux_system_env_D.master[340].sequencer;
    sequencer.master_sequencer_D341 =  pf_vf_mux_system_env_D.master[341].sequencer;
    sequencer.master_sequencer_D342 =  pf_vf_mux_system_env_D.master[342].sequencer;
    sequencer.master_sequencer_D343 =  pf_vf_mux_system_env_D.master[343].sequencer;
    sequencer.master_sequencer_D344 =  pf_vf_mux_system_env_D.master[344].sequencer;
    sequencer.master_sequencer_D345 =  pf_vf_mux_system_env_D.master[345].sequencer;
    sequencer.master_sequencer_D346 =  pf_vf_mux_system_env_D.master[346].sequencer;
    sequencer.master_sequencer_D347 =  pf_vf_mux_system_env_D.master[347].sequencer;
    sequencer.master_sequencer_D348 =  pf_vf_mux_system_env_D.master[348].sequencer;
    sequencer.master_sequencer_D349 =  pf_vf_mux_system_env_D.master[349].sequencer;
    sequencer.master_sequencer_D350 =  pf_vf_mux_system_env_D.master[350].sequencer;
    sequencer.master_sequencer_D351 =  pf_vf_mux_system_env_D.master[351].sequencer;
    sequencer.master_sequencer_D352 =  pf_vf_mux_system_env_D.master[352].sequencer;
    sequencer.master_sequencer_D353 =  pf_vf_mux_system_env_D.master[353].sequencer;
    sequencer.master_sequencer_D354 =  pf_vf_mux_system_env_D.master[354].sequencer;
    sequencer.master_sequencer_D355 =  pf_vf_mux_system_env_D.master[355].sequencer;
    sequencer.master_sequencer_D356 =  pf_vf_mux_system_env_D.master[356].sequencer;
    sequencer.master_sequencer_D357 =  pf_vf_mux_system_env_D.master[357].sequencer;
    sequencer.master_sequencer_D358 =  pf_vf_mux_system_env_D.master[358].sequencer;
    sequencer.master_sequencer_D359 =  pf_vf_mux_system_env_D.master[359].sequencer;
    sequencer.master_sequencer_D360 =  pf_vf_mux_system_env_D.master[360].sequencer;
    sequencer.master_sequencer_D361 =  pf_vf_mux_system_env_D.master[361].sequencer;
    sequencer.master_sequencer_D362 =  pf_vf_mux_system_env_D.master[362].sequencer;
    sequencer.master_sequencer_D363 =  pf_vf_mux_system_env_D.master[363].sequencer;
    sequencer.master_sequencer_D364 =  pf_vf_mux_system_env_D.master[364].sequencer;
    sequencer.master_sequencer_D365 =  pf_vf_mux_system_env_D.master[365].sequencer;
    sequencer.master_sequencer_D366 =  pf_vf_mux_system_env_D.master[366].sequencer;
    sequencer.master_sequencer_D367 =  pf_vf_mux_system_env_D.master[367].sequencer;
    sequencer.master_sequencer_D368 =  pf_vf_mux_system_env_D.master[368].sequencer;
    sequencer.master_sequencer_D369 =  pf_vf_mux_system_env_D.master[369].sequencer;
    sequencer.master_sequencer_D370 =  pf_vf_mux_system_env_D.master[370].sequencer;
    sequencer.master_sequencer_D371 =  pf_vf_mux_system_env_D.master[371].sequencer;
    sequencer.master_sequencer_D372 =  pf_vf_mux_system_env_D.master[372].sequencer;
    sequencer.master_sequencer_D373 =  pf_vf_mux_system_env_D.master[373].sequencer;
    sequencer.master_sequencer_D374 =  pf_vf_mux_system_env_D.master[374].sequencer;
    sequencer.master_sequencer_D375 =  pf_vf_mux_system_env_D.master[375].sequencer;
    sequencer.master_sequencer_D376 =  pf_vf_mux_system_env_D.master[376].sequencer;
    sequencer.master_sequencer_D377 =  pf_vf_mux_system_env_D.master[377].sequencer;
    sequencer.master_sequencer_D378 =  pf_vf_mux_system_env_D.master[378].sequencer;
    sequencer.master_sequencer_D379 =  pf_vf_mux_system_env_D.master[379].sequencer;
    sequencer.master_sequencer_D380 =  pf_vf_mux_system_env_D.master[380].sequencer;
    sequencer.master_sequencer_D381 =  pf_vf_mux_system_env_D.master[381].sequencer;
    sequencer.master_sequencer_D382 =  pf_vf_mux_system_env_D.master[382].sequencer;
    sequencer.master_sequencer_D383 =  pf_vf_mux_system_env_D.master[383].sequencer;
    sequencer.master_sequencer_D384 =  pf_vf_mux_system_env_D.master[384].sequencer;
    sequencer.master_sequencer_D385 =  pf_vf_mux_system_env_D.master[385].sequencer;
    sequencer.master_sequencer_D386 =  pf_vf_mux_system_env_D.master[386].sequencer;
    sequencer.master_sequencer_D387 =  pf_vf_mux_system_env_D.master[387].sequencer;
    sequencer.master_sequencer_D388 =  pf_vf_mux_system_env_D.master[388].sequencer;
    sequencer.master_sequencer_D389 =  pf_vf_mux_system_env_D.master[389].sequencer;
    sequencer.master_sequencer_D390 =  pf_vf_mux_system_env_D.master[390].sequencer;
    sequencer.master_sequencer_D391 =  pf_vf_mux_system_env_D.master[391].sequencer;
    sequencer.master_sequencer_D392 =  pf_vf_mux_system_env_D.master[392].sequencer;
    sequencer.master_sequencer_D393 =  pf_vf_mux_system_env_D.master[393].sequencer;
    sequencer.master_sequencer_D394 =  pf_vf_mux_system_env_D.master[394].sequencer;
    sequencer.master_sequencer_D395 =  pf_vf_mux_system_env_D.master[395].sequencer;
    sequencer.master_sequencer_D396 =  pf_vf_mux_system_env_D.master[396].sequencer;
    sequencer.master_sequencer_D397 =  pf_vf_mux_system_env_D.master[397].sequencer;
    sequencer.master_sequencer_D398 =  pf_vf_mux_system_env_D.master[398].sequencer;
    sequencer.master_sequencer_D399 =  pf_vf_mux_system_env_D.master[399].sequencer;
    sequencer.master_sequencer_D400 =  pf_vf_mux_system_env_D.master[400].sequencer;
    sequencer.master_sequencer_D401 =  pf_vf_mux_system_env_D.master[401].sequencer;
    sequencer.master_sequencer_D402 =  pf_vf_mux_system_env_D.master[402].sequencer;
    sequencer.master_sequencer_D403 =  pf_vf_mux_system_env_D.master[403].sequencer;
    sequencer.master_sequencer_D404 =  pf_vf_mux_system_env_D.master[404].sequencer;
    sequencer.master_sequencer_D405 =  pf_vf_mux_system_env_D.master[405].sequencer;
    sequencer.master_sequencer_D406 =  pf_vf_mux_system_env_D.master[406].sequencer;
    sequencer.master_sequencer_D407 =  pf_vf_mux_system_env_D.master[407].sequencer;
    sequencer.master_sequencer_D408 =  pf_vf_mux_system_env_D.master[408].sequencer;
    sequencer.master_sequencer_D409 =  pf_vf_mux_system_env_D.master[409].sequencer;
    sequencer.master_sequencer_D410 =  pf_vf_mux_system_env_D.master[410].sequencer;
    sequencer.master_sequencer_D411 =  pf_vf_mux_system_env_D.master[411].sequencer;
    sequencer.master_sequencer_D412 =  pf_vf_mux_system_env_D.master[412].sequencer;
    sequencer.master_sequencer_D413 =  pf_vf_mux_system_env_D.master[413].sequencer;
    sequencer.master_sequencer_D414 =  pf_vf_mux_system_env_D.master[414].sequencer;
    sequencer.master_sequencer_D415 =  pf_vf_mux_system_env_D.master[415].sequencer;
    sequencer.master_sequencer_D416 =  pf_vf_mux_system_env_D.master[416].sequencer;
    sequencer.master_sequencer_D417 =  pf_vf_mux_system_env_D.master[417].sequencer;
    sequencer.master_sequencer_D418 =  pf_vf_mux_system_env_D.master[418].sequencer;
    sequencer.master_sequencer_D419 =  pf_vf_mux_system_env_D.master[419].sequencer;
    sequencer.master_sequencer_D420 =  pf_vf_mux_system_env_D.master[420].sequencer;
    sequencer.master_sequencer_D421 =  pf_vf_mux_system_env_D.master[421].sequencer;
    sequencer.master_sequencer_D422 =  pf_vf_mux_system_env_D.master[422].sequencer;
    sequencer.master_sequencer_D423 =  pf_vf_mux_system_env_D.master[423].sequencer;
    sequencer.master_sequencer_D424 =  pf_vf_mux_system_env_D.master[424].sequencer;
    sequencer.master_sequencer_D425 =  pf_vf_mux_system_env_D.master[425].sequencer;
    sequencer.master_sequencer_D426 =  pf_vf_mux_system_env_D.master[426].sequencer;
    sequencer.master_sequencer_D427 =  pf_vf_mux_system_env_D.master[427].sequencer;
    sequencer.master_sequencer_D428 =  pf_vf_mux_system_env_D.master[428].sequencer;
    sequencer.master_sequencer_D429 =  pf_vf_mux_system_env_D.master[429].sequencer;
    sequencer.master_sequencer_D430 =  pf_vf_mux_system_env_D.master[430].sequencer;
    sequencer.master_sequencer_D431 =  pf_vf_mux_system_env_D.master[431].sequencer;
    sequencer.master_sequencer_D432 =  pf_vf_mux_system_env_D.master[432].sequencer;
    sequencer.master_sequencer_D433 =  pf_vf_mux_system_env_D.master[433].sequencer;
    sequencer.master_sequencer_D434 =  pf_vf_mux_system_env_D.master[434].sequencer;
    sequencer.master_sequencer_D435 =  pf_vf_mux_system_env_D.master[435].sequencer;
    sequencer.master_sequencer_D436 =  pf_vf_mux_system_env_D.master[436].sequencer;
    sequencer.master_sequencer_D437 =  pf_vf_mux_system_env_D.master[437].sequencer;
    sequencer.master_sequencer_D438 =  pf_vf_mux_system_env_D.master[438].sequencer;
    sequencer.master_sequencer_D439 =  pf_vf_mux_system_env_D.master[439].sequencer;
    sequencer.master_sequencer_D440 =  pf_vf_mux_system_env_D.master[440].sequencer;
    sequencer.master_sequencer_D441 =  pf_vf_mux_system_env_D.master[441].sequencer;
    sequencer.master_sequencer_D442 =  pf_vf_mux_system_env_D.master[442].sequencer;
    sequencer.master_sequencer_D443 =  pf_vf_mux_system_env_D.master[443].sequencer;
    sequencer.master_sequencer_D444 =  pf_vf_mux_system_env_D.master[444].sequencer;
    sequencer.master_sequencer_D445 =  pf_vf_mux_system_env_D.master[445].sequencer;
    sequencer.master_sequencer_D446 =  pf_vf_mux_system_env_D.master[446].sequencer;
    sequencer.master_sequencer_D447 =  pf_vf_mux_system_env_D.master[447].sequencer;
    sequencer.master_sequencer_D448 =  pf_vf_mux_system_env_D.master[448].sequencer;
    sequencer.master_sequencer_D449 =  pf_vf_mux_system_env_D.master[449].sequencer;
    sequencer.master_sequencer_D450 =  pf_vf_mux_system_env_TB4_D0.master[0].sequencer;
    sequencer.master_sequencer_D451 =  pf_vf_mux_system_env_TB4_D0.master[1].sequencer;
    sequencer.master_sequencer_D452 =  pf_vf_mux_system_env_TB4_D0.master[2].sequencer;
    sequencer.master_sequencer_D453 =  pf_vf_mux_system_env_TB4_D0.master[3].sequencer;
    sequencer.master_sequencer_D454 =  pf_vf_mux_system_env_TB4_D0.master[4].sequencer;
    sequencer.master_sequencer_D455 =  pf_vf_mux_system_env_TB4_D0.master[5].sequencer;
    sequencer.master_sequencer_D456 =  pf_vf_mux_system_env_TB4_D0.master[6].sequencer;
    sequencer.master_sequencer_D457 =  pf_vf_mux_system_env_TB4_D0.master[7].sequencer;
    sequencer.master_sequencer_D458 =  pf_vf_mux_system_env_TB4_D0.master[8].sequencer;
    sequencer.master_sequencer_D459 =  pf_vf_mux_system_env_TB4_D0.master[9].sequencer;
    sequencer.master_sequencer_D460 =  pf_vf_mux_system_env_TB4_D0.master[10].sequencer;
    sequencer.master_sequencer_D461 =  pf_vf_mux_system_env_TB4_D0.master[11].sequencer;
    sequencer.master_sequencer_D462 =  pf_vf_mux_system_env_TB4_D0.master[12].sequencer;
    sequencer.master_sequencer_D463 =  pf_vf_mux_system_env_TB4_D0.master[13].sequencer;
    sequencer.master_sequencer_D464 =  pf_vf_mux_system_env_TB4_D0.master[14].sequencer;
    sequencer.master_sequencer_D465 =  pf_vf_mux_system_env_TB4_D0.master[15].sequencer;
    sequencer.master_sequencer_D466 =  pf_vf_mux_system_env_TB4_D0.master[16].sequencer;
    sequencer.master_sequencer_D467 =  pf_vf_mux_system_env_TB4_D0.master[17].sequencer;
    sequencer.master_sequencer_D468 =  pf_vf_mux_system_env_TB4_D0.master[18].sequencer;
    sequencer.master_sequencer_D469 =  pf_vf_mux_system_env_TB4_D0.master[19].sequencer;
    sequencer.master_sequencer_D470 =  pf_vf_mux_system_env_TB4_D0.master[20].sequencer;
    sequencer.master_sequencer_D471 =  pf_vf_mux_system_env_TB4_D0.master[21].sequencer;
    sequencer.master_sequencer_D472 =  pf_vf_mux_system_env_TB4_D0.master[22].sequencer;
    sequencer.master_sequencer_D473 =  pf_vf_mux_system_env_TB4_D0.master[23].sequencer;
    sequencer.master_sequencer_D474 =  pf_vf_mux_system_env_TB4_D0.master[24].sequencer;
    sequencer.master_sequencer_D475 =  pf_vf_mux_system_env_TB4_D0.master[25].sequencer;
    sequencer.master_sequencer_D476 =  pf_vf_mux_system_env_TB4_D0.master[26].sequencer;
    sequencer.master_sequencer_D477 =  pf_vf_mux_system_env_TB4_D0.master[27].sequencer;
    sequencer.master_sequencer_D478 =  pf_vf_mux_system_env_TB4_D0.master[28].sequencer;
    sequencer.master_sequencer_D479 =  pf_vf_mux_system_env_TB4_D0.master[29].sequencer;
    sequencer.master_sequencer_D480 =  pf_vf_mux_system_env_TB4_D0.master[30].sequencer;
    sequencer.master_sequencer_D481 =  pf_vf_mux_system_env_TB4_D0.master[31].sequencer;
    sequencer.master_sequencer_D482 =  pf_vf_mux_system_env_TB4_D0.master[32].sequencer;
    sequencer.master_sequencer_D483 =  pf_vf_mux_system_env_TB4_D0.master[33].sequencer;
    sequencer.master_sequencer_D484 =  pf_vf_mux_system_env_TB4_D0.master[34].sequencer;
    sequencer.master_sequencer_D485 =  pf_vf_mux_system_env_TB4_D0.master[35].sequencer;
    sequencer.master_sequencer_D486 =  pf_vf_mux_system_env_TB4_D0.master[36].sequencer;
    sequencer.master_sequencer_D487 =  pf_vf_mux_system_env_TB4_D0.master[37].sequencer;
    sequencer.master_sequencer_D488 =  pf_vf_mux_system_env_TB4_D0.master[38].sequencer;
    sequencer.master_sequencer_D489 =  pf_vf_mux_system_env_TB4_D0.master[39].sequencer;
    sequencer.master_sequencer_D490 =  pf_vf_mux_system_env_TB4_D0.master[40].sequencer;
    sequencer.master_sequencer_D491 =  pf_vf_mux_system_env_TB4_D0.master[41].sequencer;
    sequencer.master_sequencer_D492 =  pf_vf_mux_system_env_TB4_D0.master[42].sequencer;
    sequencer.master_sequencer_D493 =  pf_vf_mux_system_env_TB4_D0.master[43].sequencer;
    sequencer.master_sequencer_D494 =  pf_vf_mux_system_env_TB4_D0.master[44].sequencer;
    sequencer.master_sequencer_D495 =  pf_vf_mux_system_env_TB4_D0.master[45].sequencer;
    sequencer.master_sequencer_D496 =  pf_vf_mux_system_env_TB4_D0.master[46].sequencer;
    sequencer.master_sequencer_D497 =  pf_vf_mux_system_env_TB4_D0.master[47].sequencer;
    sequencer.master_sequencer_D498 =  pf_vf_mux_system_env_TB4_D0.master[48].sequencer;
    sequencer.master_sequencer_D499 =  pf_vf_mux_system_env_TB4_D0.master[49].sequencer;
    sequencer.master_sequencer_D500 =  pf_vf_mux_system_env_TB4_D0.master[50].sequencer;
    sequencer.master_sequencer_D501 =  pf_vf_mux_system_env_TB4_D0.master[51].sequencer;
    sequencer.master_sequencer_D502 =  pf_vf_mux_system_env_TB4_D0.master[52].sequencer;
    sequencer.master_sequencer_D503 =  pf_vf_mux_system_env_TB4_D0.master[53].sequencer;
    sequencer.master_sequencer_D504 =  pf_vf_mux_system_env_TB4_D0.master[54].sequencer;
    sequencer.master_sequencer_D505 =  pf_vf_mux_system_env_TB4_D0.master[55].sequencer;
    sequencer.master_sequencer_D506 =  pf_vf_mux_system_env_TB4_D0.master[56].sequencer;
    sequencer.master_sequencer_D507 =  pf_vf_mux_system_env_TB4_D0.master[57].sequencer;
    sequencer.master_sequencer_D508 =  pf_vf_mux_system_env_TB4_D0.master[58].sequencer;
    sequencer.master_sequencer_D509 =  pf_vf_mux_system_env_TB4_D0.master[59].sequencer;
    sequencer.master_sequencer_D510 =  pf_vf_mux_system_env_TB4_D0.master[60].sequencer;
    sequencer.master_sequencer_D511 =  pf_vf_mux_system_env_TB4_D0.master[61].sequencer;
    sequencer.master_sequencer_D512 =  pf_vf_mux_system_env_TB4_D0.master[62].sequencer;
    sequencer.master_sequencer_D513 =  pf_vf_mux_system_env_TB4_D0.master[63].sequencer;
    sequencer.master_sequencer_D514 =  pf_vf_mux_system_env_TB4_D0.master[64].sequencer;
    sequencer.master_sequencer_D515 =  pf_vf_mux_system_env_TB4_D0.master[65].sequencer;
    sequencer.master_sequencer_D516 =  pf_vf_mux_system_env_TB4_D0.master[66].sequencer;
    sequencer.master_sequencer_D517 =  pf_vf_mux_system_env_TB4_D0.master[67].sequencer;
    sequencer.master_sequencer_D518 =  pf_vf_mux_system_env_TB4_D0.master[68].sequencer;
    sequencer.master_sequencer_D519 =  pf_vf_mux_system_env_TB4_D0.master[69].sequencer;
    sequencer.master_sequencer_D520 =  pf_vf_mux_system_env_TB4_D0.master[70].sequencer;
    sequencer.master_sequencer_D521 =  pf_vf_mux_system_env_TB4_D0.master[71].sequencer;
    sequencer.master_sequencer_D522 =  pf_vf_mux_system_env_TB4_D0.master[72].sequencer;
    sequencer.master_sequencer_D523 =  pf_vf_mux_system_env_TB4_D0.master[73].sequencer;
    sequencer.master_sequencer_D524 =  pf_vf_mux_system_env_TB4_D0.master[74].sequencer;
    sequencer.master_sequencer_D525 =  pf_vf_mux_system_env_TB4_D0.master[75].sequencer;
    sequencer.master_sequencer_D526 =  pf_vf_mux_system_env_TB4_D0.master[76].sequencer;
    sequencer.master_sequencer_D527 =  pf_vf_mux_system_env_TB4_D0.master[77].sequencer;
    sequencer.master_sequencer_D528 =  pf_vf_mux_system_env_TB4_D0.master[78].sequencer;
    sequencer.master_sequencer_D529 =  pf_vf_mux_system_env_TB4_D0.master[79].sequencer;
    sequencer.master_sequencer_D530 =  pf_vf_mux_system_env_TB4_D0.master[80].sequencer;
    sequencer.master_sequencer_D531 =  pf_vf_mux_system_env_TB4_D0.master[81].sequencer;
    sequencer.master_sequencer_D532 =  pf_vf_mux_system_env_TB4_D0.master[82].sequencer;
    sequencer.master_sequencer_D533 =  pf_vf_mux_system_env_TB4_D0.master[83].sequencer;
    sequencer.master_sequencer_D534 =  pf_vf_mux_system_env_TB4_D0.master[84].sequencer;
    sequencer.master_sequencer_D535 =  pf_vf_mux_system_env_TB4_D0.master[85].sequencer;
    sequencer.master_sequencer_D536 =  pf_vf_mux_system_env_TB4_D0.master[86].sequencer;
    sequencer.master_sequencer_D537 =  pf_vf_mux_system_env_TB4_D0.master[87].sequencer;
    sequencer.master_sequencer_D538 =  pf_vf_mux_system_env_TB4_D0.master[88].sequencer;
    sequencer.master_sequencer_D539 =  pf_vf_mux_system_env_TB4_D0.master[89].sequencer;
    sequencer.master_sequencer_D540 =  pf_vf_mux_system_env_TB4_D0.master[90].sequencer;
    sequencer.master_sequencer_D541 =  pf_vf_mux_system_env_TB4_D0.master[91].sequencer;
    sequencer.master_sequencer_D542 =  pf_vf_mux_system_env_TB4_D0.master[92].sequencer;
    sequencer.master_sequencer_D543 =  pf_vf_mux_system_env_TB4_D0.master[93].sequencer;
    sequencer.master_sequencer_D544 =  pf_vf_mux_system_env_TB4_D0.master[94].sequencer;
    sequencer.master_sequencer_D545 =  pf_vf_mux_system_env_TB4_D0.master[95].sequencer;
    sequencer.master_sequencer_D546 =  pf_vf_mux_system_env_TB4_D0.master[96].sequencer;
    sequencer.master_sequencer_D547 =  pf_vf_mux_system_env_TB4_D0.master[97].sequencer;
    sequencer.master_sequencer_D548 =  pf_vf_mux_system_env_TB4_D0.master[98].sequencer;
    sequencer.master_sequencer_D549 =  pf_vf_mux_system_env_TB4_D0.master[99].sequencer;
    sequencer.master_sequencer_D550 =  pf_vf_mux_system_env_TB4_D0.master[100].sequencer;
    sequencer.master_sequencer_D551 =  pf_vf_mux_system_env_TB4_D0.master[101].sequencer;
    sequencer.master_sequencer_D552 =  pf_vf_mux_system_env_TB4_D0.master[102].sequencer;
    sequencer.master_sequencer_D553 =  pf_vf_mux_system_env_TB4_D0.master[103].sequencer;
    sequencer.master_sequencer_D554 =  pf_vf_mux_system_env_TB4_D0.master[104].sequencer;
    sequencer.master_sequencer_D555 =  pf_vf_mux_system_env_TB4_D0.master[105].sequencer;
    sequencer.master_sequencer_D556 =  pf_vf_mux_system_env_TB4_D0.master[106].sequencer;
    sequencer.master_sequencer_D557 =  pf_vf_mux_system_env_TB4_D0.master[107].sequencer;
    sequencer.master_sequencer_D558 =  pf_vf_mux_system_env_TB4_D0.master[108].sequencer;
    sequencer.master_sequencer_D559 =  pf_vf_mux_system_env_TB4_D0.master[109].sequencer;
    sequencer.master_sequencer_D560 =  pf_vf_mux_system_env_TB4_D0.master[110].sequencer;
    sequencer.master_sequencer_D561 =  pf_vf_mux_system_env_TB4_D0.master[111].sequencer;
    sequencer.master_sequencer_D562 =  pf_vf_mux_system_env_TB4_D0.master[112].sequencer;
    sequencer.master_sequencer_D563 =  pf_vf_mux_system_env_TB4_D0.master[113].sequencer;
    sequencer.master_sequencer_D564 =  pf_vf_mux_system_env_TB4_D0.master[114].sequencer;
    sequencer.master_sequencer_D565 =  pf_vf_mux_system_env_TB4_D0.master[115].sequencer;
    sequencer.master_sequencer_D566 =  pf_vf_mux_system_env_TB4_D0.master[116].sequencer;
    sequencer.master_sequencer_D567 =  pf_vf_mux_system_env_TB4_D0.master[117].sequencer;
    sequencer.master_sequencer_D568 =  pf_vf_mux_system_env_TB4_D0.master[118].sequencer;
    sequencer.master_sequencer_D569 =  pf_vf_mux_system_env_TB4_D0.master[119].sequencer;
    sequencer.master_sequencer_D570 =  pf_vf_mux_system_env_TB4_D0.master[120].sequencer;
    sequencer.master_sequencer_D571 =  pf_vf_mux_system_env_TB4_D0.master[121].sequencer;
    sequencer.master_sequencer_D572 =  pf_vf_mux_system_env_TB4_D0.master[122].sequencer;
    sequencer.master_sequencer_D573 =  pf_vf_mux_system_env_TB4_D0.master[123].sequencer;
    sequencer.master_sequencer_D574 =  pf_vf_mux_system_env_TB4_D0.master[124].sequencer;
    sequencer.master_sequencer_D575 =  pf_vf_mux_system_env_TB4_D0.master[125].sequencer;
    sequencer.master_sequencer_D576 =  pf_vf_mux_system_env_TB4_D0.master[126].sequencer;
    sequencer.master_sequencer_D577 =  pf_vf_mux_system_env_TB4_D0.master[127].sequencer;
    sequencer.master_sequencer_D578 =  pf_vf_mux_system_env_TB4_D0.master[128].sequencer;
    sequencer.master_sequencer_D579 =  pf_vf_mux_system_env_TB4_D0.master[129].sequencer;
    sequencer.master_sequencer_D580 =  pf_vf_mux_system_env_TB4_D0.master[130].sequencer;
    sequencer.master_sequencer_D581 =  pf_vf_mux_system_env_TB4_D0.master[131].sequencer;
    sequencer.master_sequencer_D582 =  pf_vf_mux_system_env_TB4_D0.master[132].sequencer;
    sequencer.master_sequencer_D583 =  pf_vf_mux_system_env_TB4_D0.master[133].sequencer;
    sequencer.master_sequencer_D584 =  pf_vf_mux_system_env_TB4_D0.master[134].sequencer;
    sequencer.master_sequencer_D585 =  pf_vf_mux_system_env_TB4_D0.master[135].sequencer;
    sequencer.master_sequencer_D586 =  pf_vf_mux_system_env_TB4_D0.master[136].sequencer;
    sequencer.master_sequencer_D587 =  pf_vf_mux_system_env_TB4_D0.master[137].sequencer;
    sequencer.master_sequencer_D588 =  pf_vf_mux_system_env_TB4_D0.master[138].sequencer;
    sequencer.master_sequencer_D589 =  pf_vf_mux_system_env_TB4_D0.master[139].sequencer;
    sequencer.master_sequencer_D590 =  pf_vf_mux_system_env_TB4_D0.master[140].sequencer;
    sequencer.master_sequencer_D591 =  pf_vf_mux_system_env_TB4_D0.master[141].sequencer;
    sequencer.master_sequencer_D592 =  pf_vf_mux_system_env_TB4_D0.master[142].sequencer;
    sequencer.master_sequencer_D593 =  pf_vf_mux_system_env_TB4_D0.master[143].sequencer;
    sequencer.master_sequencer_D594 =  pf_vf_mux_system_env_TB4_D0.master[144].sequencer;
    sequencer.master_sequencer_D595 =  pf_vf_mux_system_env_TB4_D0.master[145].sequencer;
    sequencer.master_sequencer_D596 =  pf_vf_mux_system_env_TB4_D0.master[146].sequencer;
    sequencer.master_sequencer_D597 =  pf_vf_mux_system_env_TB4_D0.master[147].sequencer;
    sequencer.master_sequencer_D598 =  pf_vf_mux_system_env_TB4_D0.master[148].sequencer;
    sequencer.master_sequencer_D599 =  pf_vf_mux_system_env_TB4_D0.master[149].sequencer;
    sequencer.master_sequencer_D600 =  pf_vf_mux_system_env_TB4_D0.master[150].sequencer;
    sequencer.master_sequencer_D601 =  pf_vf_mux_system_env_TB4_D0.master[151].sequencer;
    sequencer.master_sequencer_D602 =  pf_vf_mux_system_env_TB4_D0.master[152].sequencer;
    sequencer.master_sequencer_D603 =  pf_vf_mux_system_env_TB4_D0.master[153].sequencer;
    sequencer.master_sequencer_D604 =  pf_vf_mux_system_env_TB4_D0.master[154].sequencer;
    sequencer.master_sequencer_D605 =  pf_vf_mux_system_env_TB4_D0.master[155].sequencer;
    sequencer.master_sequencer_D606 =  pf_vf_mux_system_env_TB4_D0.master[156].sequencer;
    sequencer.master_sequencer_D607 =  pf_vf_mux_system_env_TB4_D0.master[157].sequencer;
    sequencer.master_sequencer_D608 =  pf_vf_mux_system_env_TB4_D0.master[158].sequencer;
    sequencer.master_sequencer_D609 =  pf_vf_mux_system_env_TB4_D0.master[159].sequencer;
    sequencer.master_sequencer_D610 =  pf_vf_mux_system_env_TB4_D0.master[160].sequencer;
    sequencer.master_sequencer_D611 =  pf_vf_mux_system_env_TB4_D0.master[161].sequencer;
    sequencer.master_sequencer_D612 =  pf_vf_mux_system_env_TB4_D0.master[162].sequencer;
    sequencer.master_sequencer_D613 =  pf_vf_mux_system_env_TB4_D0.master[163].sequencer;
    sequencer.master_sequencer_D614 =  pf_vf_mux_system_env_TB4_D0.master[164].sequencer;
    sequencer.master_sequencer_D615 =  pf_vf_mux_system_env_TB4_D0.master[165].sequencer;
    sequencer.master_sequencer_D616 =  pf_vf_mux_system_env_TB4_D0.master[166].sequencer;
    sequencer.master_sequencer_D617 =  pf_vf_mux_system_env_TB4_D0.master[167].sequencer;
    sequencer.master_sequencer_D618 =  pf_vf_mux_system_env_TB4_D0.master[168].sequencer;
    sequencer.master_sequencer_D619 =  pf_vf_mux_system_env_TB4_D0.master[169].sequencer;
    sequencer.master_sequencer_D620 =  pf_vf_mux_system_env_TB4_D0.master[170].sequencer;
    sequencer.master_sequencer_D621 =  pf_vf_mux_system_env_TB4_D0.master[171].sequencer;
    sequencer.master_sequencer_D622 =  pf_vf_mux_system_env_TB4_D0.master[172].sequencer;
    sequencer.master_sequencer_D623 =  pf_vf_mux_system_env_TB4_D0.master[173].sequencer;
    sequencer.master_sequencer_D624 =  pf_vf_mux_system_env_TB4_D0.master[174].sequencer;
    sequencer.master_sequencer_D625 =  pf_vf_mux_system_env_TB4_D0.master[175].sequencer;
    sequencer.master_sequencer_D626 =  pf_vf_mux_system_env_TB4_D0.master[176].sequencer;
    sequencer.master_sequencer_D627 =  pf_vf_mux_system_env_TB4_D0.master[177].sequencer;
    sequencer.master_sequencer_D628 =  pf_vf_mux_system_env_TB4_D0.master[178].sequencer;
    sequencer.master_sequencer_D629 =  pf_vf_mux_system_env_TB4_D0.master[179].sequencer;
    sequencer.master_sequencer_D630 =  pf_vf_mux_system_env_TB4_D0.master[180].sequencer;
    sequencer.master_sequencer_D631 =  pf_vf_mux_system_env_TB4_D0.master[181].sequencer;
    sequencer.master_sequencer_D632 =  pf_vf_mux_system_env_TB4_D0.master[182].sequencer;
    sequencer.master_sequencer_D633 =  pf_vf_mux_system_env_TB4_D0.master[183].sequencer;
    sequencer.master_sequencer_D634 =  pf_vf_mux_system_env_TB4_D0.master[184].sequencer;
    sequencer.master_sequencer_D635 =  pf_vf_mux_system_env_TB4_D0.master[185].sequencer;
    sequencer.master_sequencer_D636 =  pf_vf_mux_system_env_TB4_D0.master[186].sequencer;
    sequencer.master_sequencer_D637 =  pf_vf_mux_system_env_TB4_D0.master[187].sequencer;
    sequencer.master_sequencer_D638 =  pf_vf_mux_system_env_TB4_D0.master[188].sequencer;
    sequencer.master_sequencer_D639 =  pf_vf_mux_system_env_TB4_D0.master[189].sequencer;
    sequencer.master_sequencer_D640 =  pf_vf_mux_system_env_TB4_D0.master[190].sequencer;
    sequencer.master_sequencer_D641 =  pf_vf_mux_system_env_TB4_D0.master[191].sequencer;
    sequencer.master_sequencer_D642 =  pf_vf_mux_system_env_TB4_D0.master[192].sequencer;
    sequencer.master_sequencer_D643 =  pf_vf_mux_system_env_TB4_D0.master[193].sequencer;
    sequencer.master_sequencer_D644 =  pf_vf_mux_system_env_TB4_D0.master[194].sequencer;
    sequencer.master_sequencer_D645 =  pf_vf_mux_system_env_TB4_D0.master[195].sequencer;
    sequencer.master_sequencer_D646 =  pf_vf_mux_system_env_TB4_D0.master[196].sequencer;
    sequencer.master_sequencer_D647 =  pf_vf_mux_system_env_TB4_D0.master[197].sequencer;
    sequencer.master_sequencer_D648 =  pf_vf_mux_system_env_TB4_D0.master[198].sequencer;
    sequencer.master_sequencer_D649 =  pf_vf_mux_system_env_TB4_D0.master[199].sequencer;
    sequencer.master_sequencer_D650 =  pf_vf_mux_system_env_TB4_D0.master[200].sequencer;
    sequencer.master_sequencer_D651 =  pf_vf_mux_system_env_TB4_D0.master[201].sequencer;
    sequencer.master_sequencer_D652 =  pf_vf_mux_system_env_TB4_D0.master[202].sequencer;
    sequencer.master_sequencer_D653 =  pf_vf_mux_system_env_TB4_D0.master[203].sequencer;
    sequencer.master_sequencer_D654 =  pf_vf_mux_system_env_TB4_D0.master[204].sequencer;
    sequencer.master_sequencer_D655 =  pf_vf_mux_system_env_TB4_D0.master[205].sequencer;
    sequencer.master_sequencer_D656 =  pf_vf_mux_system_env_TB4_D0.master[206].sequencer;
    sequencer.master_sequencer_D657 =  pf_vf_mux_system_env_TB4_D0.master[207].sequencer;
    sequencer.master_sequencer_D658 =  pf_vf_mux_system_env_TB4_D0.master[208].sequencer;
    sequencer.master_sequencer_D659 =  pf_vf_mux_system_env_TB4_D0.master[209].sequencer;
    sequencer.master_sequencer_D660 =  pf_vf_mux_system_env_TB4_D0.master[210].sequencer;
    sequencer.master_sequencer_D661 =  pf_vf_mux_system_env_TB4_D0.master[211].sequencer;
    sequencer.master_sequencer_D662 =  pf_vf_mux_system_env_TB4_D0.master[212].sequencer;
    sequencer.master_sequencer_D663 =  pf_vf_mux_system_env_TB4_D0.master[213].sequencer;
    sequencer.master_sequencer_D664 =  pf_vf_mux_system_env_TB4_D0.master[214].sequencer;
    sequencer.master_sequencer_D665 =  pf_vf_mux_system_env_TB4_D0.master[215].sequencer;
    sequencer.master_sequencer_D666 =  pf_vf_mux_system_env_TB4_D0.master[216].sequencer;
    sequencer.master_sequencer_D667 =  pf_vf_mux_system_env_TB4_D0.master[217].sequencer;
    sequencer.master_sequencer_D668 =  pf_vf_mux_system_env_TB4_D0.master[218].sequencer;
    sequencer.master_sequencer_D669 =  pf_vf_mux_system_env_TB4_D0.master[219].sequencer;
    sequencer.master_sequencer_D670 =  pf_vf_mux_system_env_TB4_D0.master[220].sequencer;
    sequencer.master_sequencer_D671 =  pf_vf_mux_system_env_TB4_D0.master[221].sequencer;
    sequencer.master_sequencer_D672 =  pf_vf_mux_system_env_TB4_D0.master[222].sequencer;
    sequencer.master_sequencer_D673 =  pf_vf_mux_system_env_TB4_D0.master[223].sequencer;
    sequencer.master_sequencer_D674 =  pf_vf_mux_system_env_TB4_D0.master[224].sequencer;
    sequencer.master_sequencer_D675 =  pf_vf_mux_system_env_TB4_D0.master[225].sequencer;
    sequencer.master_sequencer_D676 =  pf_vf_mux_system_env_TB4_D0.master[226].sequencer;
    sequencer.master_sequencer_D677 =  pf_vf_mux_system_env_TB4_D0.master[227].sequencer;
    sequencer.master_sequencer_D678 =  pf_vf_mux_system_env_TB4_D0.master[228].sequencer;
    sequencer.master_sequencer_D679 =  pf_vf_mux_system_env_TB4_D0.master[229].sequencer;
    sequencer.master_sequencer_D680 =  pf_vf_mux_system_env_TB4_D0.master[230].sequencer;
    sequencer.master_sequencer_D681 =  pf_vf_mux_system_env_TB4_D0.master[231].sequencer;
    sequencer.master_sequencer_D682 =  pf_vf_mux_system_env_TB4_D0.master[232].sequencer;
    sequencer.master_sequencer_D683 =  pf_vf_mux_system_env_TB4_D0.master[233].sequencer;
    sequencer.master_sequencer_D684 =  pf_vf_mux_system_env_TB4_D0.master[234].sequencer;
    sequencer.master_sequencer_D685 =  pf_vf_mux_system_env_TB4_D0.master[235].sequencer;
    sequencer.master_sequencer_D686 =  pf_vf_mux_system_env_TB4_D0.master[236].sequencer;
    sequencer.master_sequencer_D687 =  pf_vf_mux_system_env_TB4_D0.master[237].sequencer;
    sequencer.master_sequencer_D688 =  pf_vf_mux_system_env_TB4_D0.master[238].sequencer;
    sequencer.master_sequencer_D689 =  pf_vf_mux_system_env_TB4_D0.master[239].sequencer;
    sequencer.master_sequencer_D690 =  pf_vf_mux_system_env_TB4_D0.master[240].sequencer;
    sequencer.master_sequencer_D691 =  pf_vf_mux_system_env_TB4_D0.master[241].sequencer;
    sequencer.master_sequencer_D692 =  pf_vf_mux_system_env_TB4_D0.master[242].sequencer;
    sequencer.master_sequencer_D693 =  pf_vf_mux_system_env_TB4_D0.master[243].sequencer;
    sequencer.master_sequencer_D694 =  pf_vf_mux_system_env_TB4_D0.master[244].sequencer;
    sequencer.master_sequencer_D695 =  pf_vf_mux_system_env_TB4_D0.master[245].sequencer;
    sequencer.master_sequencer_D696 =  pf_vf_mux_system_env_TB4_D0.master[246].sequencer;
    sequencer.master_sequencer_D697 =  pf_vf_mux_system_env_TB4_D0.master[247].sequencer;
    sequencer.master_sequencer_D698 =  pf_vf_mux_system_env_TB4_D0.master[248].sequencer;
    sequencer.master_sequencer_D699 =  pf_vf_mux_system_env_TB4_D0.master[249].sequencer;
    sequencer.master_sequencer_D700 =  pf_vf_mux_system_env_TB4_D0.master[250].sequencer;
    sequencer.master_sequencer_D701 =  pf_vf_mux_system_env_TB4_D0.master[251].sequencer;
    sequencer.master_sequencer_D702 =  pf_vf_mux_system_env_TB4_D0.master[252].sequencer;
    sequencer.master_sequencer_D703 =  pf_vf_mux_system_env_TB4_D0.master[253].sequencer;
    sequencer.master_sequencer_D704 =  pf_vf_mux_system_env_TB4_D0.master[254].sequencer;
    sequencer.master_sequencer_D705 =  pf_vf_mux_system_env_TB4_D0.master[255].sequencer;
    sequencer.master_sequencer_D706 =  pf_vf_mux_system_env_TB4_D0.master[256].sequencer;
    sequencer.master_sequencer_D707 =  pf_vf_mux_system_env_TB4_D0.master[257].sequencer;
    sequencer.master_sequencer_D708 =  pf_vf_mux_system_env_TB4_D0.master[258].sequencer;
    sequencer.master_sequencer_D709 =  pf_vf_mux_system_env_TB4_D0.master[259].sequencer;
    sequencer.master_sequencer_D710 =  pf_vf_mux_system_env_TB4_D0.master[260].sequencer;
    sequencer.master_sequencer_D711 =  pf_vf_mux_system_env_TB4_D0.master[261].sequencer;
    sequencer.master_sequencer_D712 =  pf_vf_mux_system_env_TB4_D0.master[262].sequencer;
    sequencer.master_sequencer_D713 =  pf_vf_mux_system_env_TB4_D0.master[263].sequencer;
    sequencer.master_sequencer_D714 =  pf_vf_mux_system_env_TB4_D0.master[264].sequencer;
    sequencer.master_sequencer_D715 =  pf_vf_mux_system_env_TB4_D0.master[265].sequencer;
    sequencer.master_sequencer_D716 =  pf_vf_mux_system_env_TB4_D0.master[266].sequencer;
    sequencer.master_sequencer_D717 =  pf_vf_mux_system_env_TB4_D0.master[267].sequencer;
    sequencer.master_sequencer_D718 =  pf_vf_mux_system_env_TB4_D0.master[268].sequencer;
    sequencer.master_sequencer_D719 =  pf_vf_mux_system_env_TB4_D0.master[269].sequencer;
    sequencer.master_sequencer_D720 =  pf_vf_mux_system_env_TB4_D0.master[270].sequencer;
    sequencer.master_sequencer_D721 =  pf_vf_mux_system_env_TB4_D0.master[271].sequencer;
    sequencer.master_sequencer_D722 =  pf_vf_mux_system_env_TB4_D0.master[272].sequencer;
    sequencer.master_sequencer_D723 =  pf_vf_mux_system_env_TB4_D0.master[273].sequencer;
    sequencer.master_sequencer_D724 =  pf_vf_mux_system_env_TB4_D0.master[274].sequencer;
    sequencer.master_sequencer_D725 =  pf_vf_mux_system_env_TB4_D0.master[275].sequencer;
    sequencer.master_sequencer_D726 =  pf_vf_mux_system_env_TB4_D0.master[276].sequencer;
    sequencer.master_sequencer_D727 =  pf_vf_mux_system_env_TB4_D0.master[277].sequencer;
    sequencer.master_sequencer_D728 =  pf_vf_mux_system_env_TB4_D0.master[278].sequencer;
    sequencer.master_sequencer_D729 =  pf_vf_mux_system_env_TB4_D0.master[279].sequencer;
    sequencer.master_sequencer_D730 =  pf_vf_mux_system_env_TB4_D0.master[280].sequencer;
    sequencer.master_sequencer_D731 =  pf_vf_mux_system_env_TB4_D0.master[281].sequencer;
    sequencer.master_sequencer_D732 =  pf_vf_mux_system_env_TB4_D0.master[282].sequencer;
    sequencer.master_sequencer_D733 =  pf_vf_mux_system_env_TB4_D0.master[283].sequencer;
    sequencer.master_sequencer_D734 =  pf_vf_mux_system_env_TB4_D0.master[284].sequencer;
    sequencer.master_sequencer_D735 =  pf_vf_mux_system_env_TB4_D0.master[285].sequencer;
    sequencer.master_sequencer_D736 =  pf_vf_mux_system_env_TB4_D0.master[286].sequencer;
    sequencer.master_sequencer_D737 =  pf_vf_mux_system_env_TB4_D0.master[287].sequencer;
    sequencer.master_sequencer_D738 =  pf_vf_mux_system_env_TB4_D0.master[288].sequencer;
    sequencer.master_sequencer_D739 =  pf_vf_mux_system_env_TB4_D0.master[289].sequencer;
    sequencer.master_sequencer_D740 =  pf_vf_mux_system_env_TB4_D0.master[290].sequencer;
    sequencer.master_sequencer_D741 =  pf_vf_mux_system_env_TB4_D0.master[291].sequencer;
    sequencer.master_sequencer_D742 =  pf_vf_mux_system_env_TB4_D0.master[292].sequencer;
    sequencer.master_sequencer_D743 =  pf_vf_mux_system_env_TB4_D0.master[293].sequencer;
    sequencer.master_sequencer_D744 =  pf_vf_mux_system_env_TB4_D0.master[294].sequencer;
    sequencer.master_sequencer_D745 =  pf_vf_mux_system_env_TB4_D0.master[295].sequencer;
    sequencer.master_sequencer_D746 =  pf_vf_mux_system_env_TB4_D0.master[296].sequencer;
    sequencer.master_sequencer_D747 =  pf_vf_mux_system_env_TB4_D0.master[297].sequencer;
    sequencer.master_sequencer_D748 =  pf_vf_mux_system_env_TB4_D0.master[298].sequencer;
    sequencer.master_sequencer_D749 =  pf_vf_mux_system_env_TB4_D0.master[299].sequencer;
    sequencer.master_sequencer_D750 =  pf_vf_mux_system_env_TB4_D0.master[300].sequencer;
    sequencer.master_sequencer_D751 =  pf_vf_mux_system_env_TB4_D0.master[301].sequencer;
    sequencer.master_sequencer_D752 =  pf_vf_mux_system_env_TB4_D0.master[302].sequencer;
    sequencer.master_sequencer_D753 =  pf_vf_mux_system_env_TB4_D0.master[303].sequencer;
    sequencer.master_sequencer_D754 =  pf_vf_mux_system_env_TB4_D0.master[304].sequencer;
    sequencer.master_sequencer_D755 =  pf_vf_mux_system_env_TB4_D0.master[305].sequencer;
    sequencer.master_sequencer_D756 =  pf_vf_mux_system_env_TB4_D0.master[306].sequencer;
    sequencer.master_sequencer_D757 =  pf_vf_mux_system_env_TB4_D0.master[307].sequencer;
    sequencer.master_sequencer_D758 =  pf_vf_mux_system_env_TB4_D0.master[308].sequencer;
    sequencer.master_sequencer_D759 =  pf_vf_mux_system_env_TB4_D0.master[309].sequencer;
    sequencer.master_sequencer_D760 =  pf_vf_mux_system_env_TB4_D0.master[310].sequencer;
    sequencer.master_sequencer_D761 =  pf_vf_mux_system_env_TB4_D0.master[311].sequencer;
    sequencer.master_sequencer_D762 =  pf_vf_mux_system_env_TB4_D0.master[312].sequencer;
    sequencer.master_sequencer_D763 =  pf_vf_mux_system_env_TB4_D0.master[313].sequencer;
    sequencer.master_sequencer_D764 =  pf_vf_mux_system_env_TB4_D0.master[314].sequencer;
    sequencer.master_sequencer_D765 =  pf_vf_mux_system_env_TB4_D0.master[315].sequencer;
    sequencer.master_sequencer_D766 =  pf_vf_mux_system_env_TB4_D0.master[316].sequencer;
    sequencer.master_sequencer_D767 =  pf_vf_mux_system_env_TB4_D0.master[317].sequencer;
    sequencer.master_sequencer_D768 =  pf_vf_mux_system_env_TB4_D0.master[318].sequencer;
    sequencer.master_sequencer_D769 =  pf_vf_mux_system_env_TB4_D0.master[319].sequencer;
    sequencer.master_sequencer_D770 =  pf_vf_mux_system_env_TB4_D0.master[320].sequencer;
    sequencer.master_sequencer_D771 =  pf_vf_mux_system_env_TB4_D0.master[321].sequencer;
    sequencer.master_sequencer_D772 =  pf_vf_mux_system_env_TB4_D0.master[322].sequencer;
    sequencer.master_sequencer_D773 =  pf_vf_mux_system_env_TB4_D0.master[323].sequencer;
    sequencer.master_sequencer_D774 =  pf_vf_mux_system_env_TB4_D0.master[324].sequencer;
    sequencer.master_sequencer_D775 =  pf_vf_mux_system_env_TB4_D0.master[325].sequencer;
    sequencer.master_sequencer_D776 =  pf_vf_mux_system_env_TB4_D0.master[326].sequencer;
    sequencer.master_sequencer_D777 =  pf_vf_mux_system_env_TB4_D0.master[327].sequencer;
    sequencer.master_sequencer_D778 =  pf_vf_mux_system_env_TB4_D0.master[328].sequencer;
    sequencer.master_sequencer_D779 =  pf_vf_mux_system_env_TB4_D0.master[329].sequencer;
    sequencer.master_sequencer_D780 =  pf_vf_mux_system_env_TB4_D0.master[330].sequencer;
    sequencer.master_sequencer_D781 =  pf_vf_mux_system_env_TB4_D0.master[331].sequencer;
    sequencer.master_sequencer_D782 =  pf_vf_mux_system_env_TB4_D0.master[332].sequencer;
    sequencer.master_sequencer_D783 =  pf_vf_mux_system_env_TB4_D0.master[333].sequencer;
    sequencer.master_sequencer_D784 =  pf_vf_mux_system_env_TB4_D0.master[334].sequencer;
    sequencer.master_sequencer_D785 =  pf_vf_mux_system_env_TB4_D0.master[335].sequencer;
    sequencer.master_sequencer_D786 =  pf_vf_mux_system_env_TB4_D0.master[336].sequencer;
    sequencer.master_sequencer_D787 =  pf_vf_mux_system_env_TB4_D0.master[337].sequencer;
    sequencer.master_sequencer_D788 =  pf_vf_mux_system_env_TB4_D0.master[338].sequencer;
    sequencer.master_sequencer_D789 =  pf_vf_mux_system_env_TB4_D0.master[339].sequencer;
    sequencer.master_sequencer_D790 =  pf_vf_mux_system_env_TB4_D0.master[340].sequencer;
    sequencer.master_sequencer_D791 =  pf_vf_mux_system_env_TB4_D0.master[341].sequencer;
    sequencer.master_sequencer_D792 =  pf_vf_mux_system_env_TB4_D0.master[342].sequencer;
    sequencer.master_sequencer_D793 =  pf_vf_mux_system_env_TB4_D0.master[343].sequencer;
    sequencer.master_sequencer_D794 =  pf_vf_mux_system_env_TB4_D0.master[344].sequencer;
    sequencer.master_sequencer_D795 =  pf_vf_mux_system_env_TB4_D0.master[345].sequencer;
    sequencer.master_sequencer_D796 =  pf_vf_mux_system_env_TB4_D0.master[346].sequencer;
    sequencer.master_sequencer_D797 =  pf_vf_mux_system_env_TB4_D0.master[347].sequencer;
    sequencer.master_sequencer_D798 =  pf_vf_mux_system_env_TB4_D0.master[348].sequencer;
    sequencer.master_sequencer_D799 =  pf_vf_mux_system_env_TB4_D0.master[349].sequencer;
    sequencer.master_sequencer_D800 =  pf_vf_mux_system_env_TB4_D0.master[350].sequencer;
    sequencer.master_sequencer_D801 =  pf_vf_mux_system_env_TB4_D0.master[351].sequencer;
    sequencer.master_sequencer_D802 =  pf_vf_mux_system_env_TB4_D0.master[352].sequencer;
    sequencer.master_sequencer_D803 =  pf_vf_mux_system_env_TB4_D0.master[353].sequencer;
    sequencer.master_sequencer_D804 =  pf_vf_mux_system_env_TB4_D0.master[354].sequencer;
    sequencer.master_sequencer_D805 =  pf_vf_mux_system_env_TB4_D0.master[355].sequencer;
    sequencer.master_sequencer_D806 =  pf_vf_mux_system_env_TB4_D0.master[356].sequencer;
    sequencer.master_sequencer_D807 =  pf_vf_mux_system_env_TB4_D0.master[357].sequencer;
    sequencer.master_sequencer_D808 =  pf_vf_mux_system_env_TB4_D0.master[358].sequencer;
    sequencer.master_sequencer_D809 =  pf_vf_mux_system_env_TB4_D0.master[359].sequencer;
    sequencer.master_sequencer_D810 =  pf_vf_mux_system_env_TB4_D0.master[360].sequencer;
    sequencer.master_sequencer_D811 =  pf_vf_mux_system_env_TB4_D0.master[361].sequencer;
    sequencer.master_sequencer_D812 =  pf_vf_mux_system_env_TB4_D0.master[362].sequencer;
    sequencer.master_sequencer_D813 =  pf_vf_mux_system_env_TB4_D0.master[363].sequencer;
    sequencer.master_sequencer_D814 =  pf_vf_mux_system_env_TB4_D0.master[364].sequencer;
    sequencer.master_sequencer_D815 =  pf_vf_mux_system_env_TB4_D0.master[365].sequencer;
    sequencer.master_sequencer_D816 =  pf_vf_mux_system_env_TB4_D0.master[366].sequencer;
    sequencer.master_sequencer_D817 =  pf_vf_mux_system_env_TB4_D0.master[367].sequencer;
    sequencer.master_sequencer_D818 =  pf_vf_mux_system_env_TB4_D0.master[368].sequencer;
    sequencer.master_sequencer_D819 =  pf_vf_mux_system_env_TB4_D0.master[369].sequencer;
    sequencer.master_sequencer_D820 =  pf_vf_mux_system_env_TB4_D0.master[370].sequencer;
    sequencer.master_sequencer_D821 =  pf_vf_mux_system_env_TB4_D0.master[371].sequencer;
    sequencer.master_sequencer_D822 =  pf_vf_mux_system_env_TB4_D0.master[372].sequencer;
    sequencer.master_sequencer_D823 =  pf_vf_mux_system_env_TB4_D0.master[373].sequencer;
    sequencer.master_sequencer_D824 =  pf_vf_mux_system_env_TB4_D0.master[374].sequencer;
    sequencer.master_sequencer_D825 =  pf_vf_mux_system_env_TB4_D0.master[375].sequencer;
    sequencer.master_sequencer_D826 =  pf_vf_mux_system_env_TB4_D0.master[376].sequencer;
    sequencer.master_sequencer_D827 =  pf_vf_mux_system_env_TB4_D0.master[377].sequencer;
    sequencer.master_sequencer_D828 =  pf_vf_mux_system_env_TB4_D0.master[378].sequencer;
    sequencer.master_sequencer_D829 =  pf_vf_mux_system_env_TB4_D0.master[379].sequencer;
    sequencer.master_sequencer_D830 =  pf_vf_mux_system_env_TB4_D0.master[380].sequencer;
    sequencer.master_sequencer_D831 =  pf_vf_mux_system_env_TB4_D0.master[381].sequencer;
    sequencer.master_sequencer_D832 =  pf_vf_mux_system_env_TB4_D0.master[382].sequencer;
    sequencer.master_sequencer_D833 =  pf_vf_mux_system_env_TB4_D0.master[383].sequencer;
    sequencer.master_sequencer_D834 =  pf_vf_mux_system_env_TB4_D0.master[384].sequencer;
    sequencer.master_sequencer_D835 =  pf_vf_mux_system_env_TB4_D0.master[385].sequencer;
    sequencer.master_sequencer_D836 =  pf_vf_mux_system_env_TB4_D0.master[386].sequencer;
    sequencer.master_sequencer_D837 =  pf_vf_mux_system_env_TB4_D0.master[387].sequencer;
    sequencer.master_sequencer_D838 =  pf_vf_mux_system_env_TB4_D0.master[388].sequencer;
    sequencer.master_sequencer_D839 =  pf_vf_mux_system_env_TB4_D0.master[389].sequencer;
    sequencer.master_sequencer_D840 =  pf_vf_mux_system_env_TB4_D0.master[390].sequencer;
    sequencer.master_sequencer_D841 =  pf_vf_mux_system_env_TB4_D0.master[391].sequencer;
    sequencer.master_sequencer_D842 =  pf_vf_mux_system_env_TB4_D0.master[392].sequencer;
    sequencer.master_sequencer_D843 =  pf_vf_mux_system_env_TB4_D0.master[393].sequencer;
    sequencer.master_sequencer_D844 =  pf_vf_mux_system_env_TB4_D0.master[394].sequencer;
    sequencer.master_sequencer_D845 =  pf_vf_mux_system_env_TB4_D0.master[395].sequencer;
    sequencer.master_sequencer_D846 =  pf_vf_mux_system_env_TB4_D0.master[396].sequencer;
    sequencer.master_sequencer_D847 =  pf_vf_mux_system_env_TB4_D0.master[397].sequencer;
    sequencer.master_sequencer_D848 =  pf_vf_mux_system_env_TB4_D0.master[398].sequencer;
    sequencer.master_sequencer_D849 =  pf_vf_mux_system_env_TB4_D0.master[399].sequencer;
    sequencer.master_sequencer_D850 =  pf_vf_mux_system_env_TB4_D0.master[400].sequencer;
    sequencer.master_sequencer_D851 =  pf_vf_mux_system_env_TB4_D0.master[401].sequencer;
    sequencer.master_sequencer_D852 =  pf_vf_mux_system_env_TB4_D0.master[402].sequencer;
    sequencer.master_sequencer_D853 =  pf_vf_mux_system_env_TB4_D0.master[403].sequencer;
    sequencer.master_sequencer_D854 =  pf_vf_mux_system_env_TB4_D0.master[404].sequencer;
    sequencer.master_sequencer_D855 =  pf_vf_mux_system_env_TB4_D0.master[405].sequencer;
    sequencer.master_sequencer_D856 =  pf_vf_mux_system_env_TB4_D0.master[406].sequencer;
    sequencer.master_sequencer_D857 =  pf_vf_mux_system_env_TB4_D0.master[407].sequencer;
    sequencer.master_sequencer_D858 =  pf_vf_mux_system_env_TB4_D0.master[408].sequencer;
    sequencer.master_sequencer_D859 =  pf_vf_mux_system_env_TB4_D0.master[409].sequencer;
    sequencer.master_sequencer_D860 =  pf_vf_mux_system_env_TB4_D0.master[410].sequencer;
    sequencer.master_sequencer_D861 =  pf_vf_mux_system_env_TB4_D0.master[411].sequencer;
    sequencer.master_sequencer_D862 =  pf_vf_mux_system_env_TB4_D0.master[412].sequencer;
    sequencer.master_sequencer_D863 =  pf_vf_mux_system_env_TB4_D0.master[413].sequencer;
    sequencer.master_sequencer_D864 =  pf_vf_mux_system_env_TB4_D0.master[414].sequencer;
    sequencer.master_sequencer_D865 =  pf_vf_mux_system_env_TB4_D0.master[415].sequencer;
    sequencer.master_sequencer_D866 =  pf_vf_mux_system_env_TB4_D0.master[416].sequencer;
    sequencer.master_sequencer_D867 =  pf_vf_mux_system_env_TB4_D0.master[417].sequencer;
    sequencer.master_sequencer_D868 =  pf_vf_mux_system_env_TB4_D0.master[418].sequencer;
    sequencer.master_sequencer_D869 =  pf_vf_mux_system_env_TB4_D0.master[419].sequencer;
    sequencer.master_sequencer_D870 =  pf_vf_mux_system_env_TB4_D0.master[420].sequencer;
    sequencer.master_sequencer_D871 =  pf_vf_mux_system_env_TB4_D0.master[421].sequencer;
    sequencer.master_sequencer_D872 =  pf_vf_mux_system_env_TB4_D0.master[422].sequencer;
    sequencer.master_sequencer_D873 =  pf_vf_mux_system_env_TB4_D0.master[423].sequencer;
    sequencer.master_sequencer_D874 =  pf_vf_mux_system_env_TB4_D0.master[424].sequencer;
    sequencer.master_sequencer_D875 =  pf_vf_mux_system_env_TB4_D0.master[425].sequencer;
    sequencer.master_sequencer_D876 =  pf_vf_mux_system_env_TB4_D0.master[426].sequencer;
    sequencer.master_sequencer_D877 =  pf_vf_mux_system_env_TB4_D0.master[427].sequencer;
    sequencer.master_sequencer_D878 =  pf_vf_mux_system_env_TB4_D0.master[428].sequencer;
    sequencer.master_sequencer_D879 =  pf_vf_mux_system_env_TB4_D0.master[429].sequencer;
    sequencer.master_sequencer_D880 =  pf_vf_mux_system_env_TB4_D0.master[430].sequencer;
    sequencer.master_sequencer_D881 =  pf_vf_mux_system_env_TB4_D0.master[431].sequencer;
    sequencer.master_sequencer_D882 =  pf_vf_mux_system_env_TB4_D0.master[432].sequencer;
    sequencer.master_sequencer_D883 =  pf_vf_mux_system_env_TB4_D0.master[433].sequencer;
    sequencer.master_sequencer_D884 =  pf_vf_mux_system_env_TB4_D0.master[434].sequencer;
    sequencer.master_sequencer_D885 =  pf_vf_mux_system_env_TB4_D0.master[435].sequencer;
    sequencer.master_sequencer_D886 =  pf_vf_mux_system_env_TB4_D0.master[436].sequencer;
    sequencer.master_sequencer_D887 =  pf_vf_mux_system_env_TB4_D0.master[437].sequencer;
    sequencer.master_sequencer_D888 =  pf_vf_mux_system_env_TB4_D0.master[438].sequencer;
    sequencer.master_sequencer_D889 =  pf_vf_mux_system_env_TB4_D0.master[439].sequencer;
    sequencer.master_sequencer_D890 =  pf_vf_mux_system_env_TB4_D0.master[440].sequencer;
    sequencer.master_sequencer_D891 =  pf_vf_mux_system_env_TB4_D0.master[441].sequencer;
    sequencer.master_sequencer_D892 =  pf_vf_mux_system_env_TB4_D0.master[442].sequencer;
    sequencer.master_sequencer_D893 =  pf_vf_mux_system_env_TB4_D0.master[443].sequencer;
    sequencer.master_sequencer_D894 =  pf_vf_mux_system_env_TB4_D0.master[444].sequencer;
    sequencer.master_sequencer_D895 =  pf_vf_mux_system_env_TB4_D0.master[445].sequencer;
    sequencer.master_sequencer_D896 =  pf_vf_mux_system_env_TB4_D0.master[446].sequencer;
    sequencer.master_sequencer_D897 =  pf_vf_mux_system_env_TB4_D0.master[447].sequencer;
    sequencer.master_sequencer_D898 =  pf_vf_mux_system_env_TB4_D0.master[448].sequencer;
    sequencer.master_sequencer_D899 =  pf_vf_mux_system_env_TB4_D0.master[449].sequencer;
    sequencer.master_sequencer_D900 =  pf_vf_mux_system_env_TB4_D1.master[0].sequencer;   
    sequencer.master_sequencer_D901 =  pf_vf_mux_system_env_TB4_D1.master[1].sequencer;   
    sequencer.master_sequencer_D902 =  pf_vf_mux_system_env_TB4_D1.master[2].sequencer;   
    sequencer.master_sequencer_D903 =  pf_vf_mux_system_env_TB4_D1.master[3].sequencer;   
    sequencer.master_sequencer_D904 =  pf_vf_mux_system_env_TB4_D1.master[4].sequencer;   
    sequencer.master_sequencer_D905 =  pf_vf_mux_system_env_TB4_D1.master[5].sequencer;   
    sequencer.master_sequencer_D906 =  pf_vf_mux_system_env_TB4_D1.master[6].sequencer;   
    sequencer.master_sequencer_D907 =  pf_vf_mux_system_env_TB4_D1.master[7].sequencer;   
    sequencer.master_sequencer_D908 =  pf_vf_mux_system_env_TB4_D1.master[8].sequencer;   
    sequencer.master_sequencer_D909 =  pf_vf_mux_system_env_TB4_D1.master[9].sequencer;   
    sequencer.master_sequencer_D910 =  pf_vf_mux_system_env_TB4_D1.master[10].sequencer;   
    sequencer.master_sequencer_D911 =  pf_vf_mux_system_env_TB4_D1.master[11].sequencer;   
    sequencer.master_sequencer_D912 =  pf_vf_mux_system_env_TB4_D1.master[12].sequencer;   
    sequencer.master_sequencer_D913 =  pf_vf_mux_system_env_TB4_D1.master[13].sequencer;   
    sequencer.master_sequencer_D914 =  pf_vf_mux_system_env_TB4_D1.master[14].sequencer;   
    sequencer.master_sequencer_D915 =  pf_vf_mux_system_env_TB4_D1.master[15].sequencer;   
    sequencer.master_sequencer_D916 =  pf_vf_mux_system_env_TB4_D1.master[16].sequencer;   
    sequencer.master_sequencer_D917 =  pf_vf_mux_system_env_TB4_D1.master[17].sequencer;   
    sequencer.master_sequencer_D918 =  pf_vf_mux_system_env_TB4_D1.master[18].sequencer;   
    sequencer.master_sequencer_D919 =  pf_vf_mux_system_env_TB4_D1.master[19].sequencer;   
    sequencer.master_sequencer_D920 =  pf_vf_mux_system_env_TB4_D1.master[20].sequencer;   
    sequencer.master_sequencer_D921 =  pf_vf_mux_system_env_TB4_D1.master[21].sequencer;   
    sequencer.master_sequencer_D922 =  pf_vf_mux_system_env_TB4_D1.master[22].sequencer;   
    sequencer.master_sequencer_D923 =  pf_vf_mux_system_env_TB4_D1.master[23].sequencer;   
    sequencer.master_sequencer_D924 =  pf_vf_mux_system_env_TB4_D1.master[24].sequencer;   
    sequencer.master_sequencer_D925 =  pf_vf_mux_system_env_TB4_D1.master[25].sequencer;   
    sequencer.master_sequencer_D926 =  pf_vf_mux_system_env_TB4_D1.master[26].sequencer;   
    sequencer.master_sequencer_D927 =  pf_vf_mux_system_env_TB4_D1.master[27].sequencer;   
    sequencer.master_sequencer_D928 =  pf_vf_mux_system_env_TB4_D1.master[28].sequencer;   
    sequencer.master_sequencer_D929 =  pf_vf_mux_system_env_TB4_D1.master[29].sequencer;   
    sequencer.master_sequencer_D930 =  pf_vf_mux_system_env_TB4_D1.master[30].sequencer;   
    sequencer.master_sequencer_D931 =  pf_vf_mux_system_env_TB4_D1.master[31].sequencer;   
    sequencer.master_sequencer_D932 =  pf_vf_mux_system_env_TB4_D1.master[32].sequencer;   
    sequencer.master_sequencer_D933 =  pf_vf_mux_system_env_TB4_D1.master[33].sequencer;   
    sequencer.master_sequencer_D934 =  pf_vf_mux_system_env_TB4_D1.master[34].sequencer;   
    sequencer.master_sequencer_D935 =  pf_vf_mux_system_env_TB4_D1.master[35].sequencer;   
    sequencer.master_sequencer_D936 =  pf_vf_mux_system_env_TB4_D1.master[36].sequencer;   
    sequencer.master_sequencer_D937 =  pf_vf_mux_system_env_TB4_D1.master[37].sequencer;   
    sequencer.master_sequencer_D938 =  pf_vf_mux_system_env_TB4_D1.master[38].sequencer;   
    sequencer.master_sequencer_D939 =  pf_vf_mux_system_env_TB4_D1.master[39].sequencer;   
    sequencer.master_sequencer_D940 =  pf_vf_mux_system_env_TB4_D1.master[40].sequencer;   
    sequencer.master_sequencer_D941 =  pf_vf_mux_system_env_TB4_D1.master[41].sequencer;   
    sequencer.master_sequencer_D942 =  pf_vf_mux_system_env_TB4_D1.master[42].sequencer;   
    sequencer.master_sequencer_D943 =  pf_vf_mux_system_env_TB4_D1.master[43].sequencer;   
    sequencer.master_sequencer_D944 =  pf_vf_mux_system_env_TB4_D1.master[44].sequencer;   
    sequencer.master_sequencer_D945 =  pf_vf_mux_system_env_TB4_D1.master[45].sequencer;   
    sequencer.master_sequencer_D946 =  pf_vf_mux_system_env_TB4_D1.master[46].sequencer;   
    sequencer.master_sequencer_D947 =  pf_vf_mux_system_env_TB4_D1.master[47].sequencer;   
    sequencer.master_sequencer_D948 =  pf_vf_mux_system_env_TB4_D1.master[48].sequencer;   
    sequencer.master_sequencer_D949 =  pf_vf_mux_system_env_TB4_D1.master[49].sequencer;   
    sequencer.master_sequencer_D950 =  pf_vf_mux_system_env_TB4_D1.master[50].sequencer;   
    sequencer.master_sequencer_D951 =  pf_vf_mux_system_env_TB4_D1.master[51].sequencer;   
    sequencer.master_sequencer_D952 =  pf_vf_mux_system_env_TB4_D1.master[52].sequencer;   
    sequencer.master_sequencer_D953 =  pf_vf_mux_system_env_TB4_D1.master[53].sequencer;   
    sequencer.master_sequencer_D954 =  pf_vf_mux_system_env_TB4_D1.master[54].sequencer;   
    sequencer.master_sequencer_D955 =  pf_vf_mux_system_env_TB4_D1.master[55].sequencer;   
    sequencer.master_sequencer_D956 =  pf_vf_mux_system_env_TB4_D1.master[56].sequencer;   
    sequencer.master_sequencer_D957 =  pf_vf_mux_system_env_TB4_D1.master[57].sequencer;   
    sequencer.master_sequencer_D958 =  pf_vf_mux_system_env_TB4_D1.master[58].sequencer;   
    sequencer.master_sequencer_D959 =  pf_vf_mux_system_env_TB4_D1.master[59].sequencer;   
    sequencer.master_sequencer_D960 =  pf_vf_mux_system_env_TB4_D1.master[60].sequencer;   
    sequencer.master_sequencer_D961 =  pf_vf_mux_system_env_TB4_D1.master[61].sequencer;   
    sequencer.master_sequencer_D962 =  pf_vf_mux_system_env_TB4_D1.master[62].sequencer;   
    sequencer.master_sequencer_D963 =  pf_vf_mux_system_env_TB4_D1.master[63].sequencer;   
    sequencer.master_sequencer_D964 =  pf_vf_mux_system_env_TB4_D1.master[64].sequencer;   
    sequencer.master_sequencer_D965 =  pf_vf_mux_system_env_TB4_D1.master[65].sequencer;   
    sequencer.master_sequencer_D966 =  pf_vf_mux_system_env_TB4_D1.master[66].sequencer;   
    sequencer.master_sequencer_D967 =  pf_vf_mux_system_env_TB4_D1.master[67].sequencer;   
    sequencer.master_sequencer_D968 =  pf_vf_mux_system_env_TB4_D1.master[68].sequencer;   
    sequencer.master_sequencer_D969 =  pf_vf_mux_system_env_TB4_D1.master[69].sequencer;   
    sequencer.master_sequencer_D970 =  pf_vf_mux_system_env_TB4_D1.master[70].sequencer;   
    sequencer.master_sequencer_D971 =  pf_vf_mux_system_env_TB4_D1.master[71].sequencer;   
    sequencer.master_sequencer_D972 =  pf_vf_mux_system_env_TB4_D1.master[72].sequencer;   
    sequencer.master_sequencer_D973 =  pf_vf_mux_system_env_TB4_D1.master[73].sequencer;   
    sequencer.master_sequencer_D974 =  pf_vf_mux_system_env_TB4_D1.master[74].sequencer;   
    sequencer.master_sequencer_D975 =  pf_vf_mux_system_env_TB4_D1.master[75].sequencer;   
    sequencer.master_sequencer_D976 =  pf_vf_mux_system_env_TB4_D1.master[76].sequencer;   
    sequencer.master_sequencer_D977 =  pf_vf_mux_system_env_TB4_D1.master[77].sequencer;   
    sequencer.master_sequencer_D978 =  pf_vf_mux_system_env_TB4_D1.master[78].sequencer;   
    sequencer.master_sequencer_D979 =  pf_vf_mux_system_env_TB4_D1.master[79].sequencer;   
    sequencer.master_sequencer_D980 =  pf_vf_mux_system_env_TB4_D1.master[80].sequencer;   
    sequencer.master_sequencer_D981 =  pf_vf_mux_system_env_TB4_D1.master[81].sequencer;   
    sequencer.master_sequencer_D982 =  pf_vf_mux_system_env_TB4_D1.master[82].sequencer;   
    sequencer.master_sequencer_D983 =  pf_vf_mux_system_env_TB4_D1.master[83].sequencer;   
    sequencer.master_sequencer_D984 =  pf_vf_mux_system_env_TB4_D1.master[84].sequencer;   
    sequencer.master_sequencer_D985 =  pf_vf_mux_system_env_TB4_D1.master[85].sequencer;   
    sequencer.master_sequencer_D986 =  pf_vf_mux_system_env_TB4_D1.master[86].sequencer;   
    sequencer.master_sequencer_D987 =  pf_vf_mux_system_env_TB4_D1.master[87].sequencer;   
    sequencer.master_sequencer_D988 =  pf_vf_mux_system_env_TB4_D1.master[88].sequencer;   
    sequencer.master_sequencer_D989 =  pf_vf_mux_system_env_TB4_D1.master[89].sequencer;   
    sequencer.master_sequencer_D990 =  pf_vf_mux_system_env_TB4_D1.master[90].sequencer;   
    sequencer.master_sequencer_D991 =  pf_vf_mux_system_env_TB4_D1.master[91].sequencer;   
    sequencer.master_sequencer_D992 =  pf_vf_mux_system_env_TB4_D1.master[92].sequencer;   
    sequencer.master_sequencer_D993 =  pf_vf_mux_system_env_TB4_D1.master[93].sequencer;   
    sequencer.master_sequencer_D994 =  pf_vf_mux_system_env_TB4_D1.master[94].sequencer;   
    sequencer.master_sequencer_D995 =  pf_vf_mux_system_env_TB4_D1.master[95].sequencer;   
    sequencer.master_sequencer_D996 =  pf_vf_mux_system_env_TB4_D1.master[96].sequencer;   
    sequencer.master_sequencer_D997 =  pf_vf_mux_system_env_TB4_D1.master[97].sequencer;   
    sequencer.master_sequencer_D998 =  pf_vf_mux_system_env_TB4_D1.master[98].sequencer;   
    sequencer.master_sequencer_D999 =  pf_vf_mux_system_env_TB4_D1.master[99].sequencer;   
    sequencer.master_sequencer_D1000 =  pf_vf_mux_system_env_TB4_D1.master[100].sequencer;   
    sequencer.master_sequencer_D1001 =  pf_vf_mux_system_env_TB4_D1.master[101].sequencer;   
    sequencer.master_sequencer_D1002 =  pf_vf_mux_system_env_TB4_D1.master[102].sequencer;   
    sequencer.master_sequencer_D1003 =  pf_vf_mux_system_env_TB4_D1.master[103].sequencer;   
    sequencer.master_sequencer_D1004 =  pf_vf_mux_system_env_TB4_D1.master[104].sequencer;   
    sequencer.master_sequencer_D1005 =  pf_vf_mux_system_env_TB4_D1.master[105].sequencer;   
    sequencer.master_sequencer_D1006 =  pf_vf_mux_system_env_TB4_D1.master[106].sequencer;   
    sequencer.master_sequencer_D1007 =  pf_vf_mux_system_env_TB4_D1.master[107].sequencer;   
    sequencer.master_sequencer_D1008 =  pf_vf_mux_system_env_TB4_D1.master[108].sequencer;   
    sequencer.master_sequencer_D1009 =  pf_vf_mux_system_env_TB4_D1.master[109].sequencer;   
    sequencer.master_sequencer_D1010 =  pf_vf_mux_system_env_TB4_D1.master[110].sequencer;   
    sequencer.master_sequencer_D1011 =  pf_vf_mux_system_env_TB4_D1.master[111].sequencer;   
    sequencer.master_sequencer_D1012 =  pf_vf_mux_system_env_TB4_D1.master[112].sequencer;   
    sequencer.master_sequencer_D1013 =  pf_vf_mux_system_env_TB4_D1.master[113].sequencer;   
    sequencer.master_sequencer_D1014 =  pf_vf_mux_system_env_TB4_D1.master[114].sequencer;   
    sequencer.master_sequencer_D1015 =  pf_vf_mux_system_env_TB4_D1.master[115].sequencer;   
    sequencer.master_sequencer_D1016 =  pf_vf_mux_system_env_TB4_D1.master[116].sequencer;   
    sequencer.master_sequencer_D1017 =  pf_vf_mux_system_env_TB4_D1.master[117].sequencer;   
    sequencer.master_sequencer_D1018 =  pf_vf_mux_system_env_TB4_D1.master[118].sequencer;   
    sequencer.master_sequencer_D1019 =  pf_vf_mux_system_env_TB4_D1.master[119].sequencer;   
    sequencer.master_sequencer_D1020 =  pf_vf_mux_system_env_TB4_D1.master[120].sequencer;   
    sequencer.master_sequencer_D1021 =  pf_vf_mux_system_env_TB4_D1.master[121].sequencer;   
    sequencer.master_sequencer_D1022 =  pf_vf_mux_system_env_TB4_D1.master[122].sequencer;   
    sequencer.master_sequencer_D1023 =  pf_vf_mux_system_env_TB4_D1.master[123].sequencer;   
    sequencer.master_sequencer_D1024 =  pf_vf_mux_system_env_TB4_D1.master[124].sequencer;   
    sequencer.master_sequencer_D1025 =  pf_vf_mux_system_env_TB4_D1.master[125].sequencer;   
    sequencer.master_sequencer_D1026 =  pf_vf_mux_system_env_TB4_D1.master[126].sequencer;   
    sequencer.master_sequencer_D1027 =  pf_vf_mux_system_env_TB4_D1.master[127].sequencer;   
    sequencer.master_sequencer_D1028 =  pf_vf_mux_system_env_TB4_D1.master[128].sequencer;   
    sequencer.master_sequencer_D1029 =  pf_vf_mux_system_env_TB4_D1.master[129].sequencer;   
    sequencer.master_sequencer_D1030 =  pf_vf_mux_system_env_TB4_D1.master[130].sequencer;   
    sequencer.master_sequencer_D1031 =  pf_vf_mux_system_env_TB4_D1.master[131].sequencer;   
    sequencer.master_sequencer_D1032 =  pf_vf_mux_system_env_TB4_D1.master[132].sequencer;   
    sequencer.master_sequencer_D1033 =  pf_vf_mux_system_env_TB4_D1.master[133].sequencer;   
    sequencer.master_sequencer_D1034 =  pf_vf_mux_system_env_TB4_D1.master[134].sequencer;   
    sequencer.master_sequencer_D1035 =  pf_vf_mux_system_env_TB4_D1.master[135].sequencer;   
    sequencer.master_sequencer_D1036 =  pf_vf_mux_system_env_TB4_D1.master[136].sequencer;   
    sequencer.master_sequencer_D1037 =  pf_vf_mux_system_env_TB4_D1.master[137].sequencer;   
    sequencer.master_sequencer_D1038 =  pf_vf_mux_system_env_TB4_D1.master[138].sequencer;   
    sequencer.master_sequencer_D1039 =  pf_vf_mux_system_env_TB4_D1.master[139].sequencer;   
    sequencer.master_sequencer_D1040 =  pf_vf_mux_system_env_TB4_D1.master[140].sequencer;   
    sequencer.master_sequencer_D1041 =  pf_vf_mux_system_env_TB4_D1.master[141].sequencer;   
    sequencer.master_sequencer_D1042 =  pf_vf_mux_system_env_TB4_D1.master[142].sequencer;   
    sequencer.master_sequencer_D1043 =  pf_vf_mux_system_env_TB4_D1.master[143].sequencer;   
    sequencer.master_sequencer_D1044 =  pf_vf_mux_system_env_TB4_D1.master[144].sequencer;   
    sequencer.master_sequencer_D1045 =  pf_vf_mux_system_env_TB4_D1.master[145].sequencer;   
    sequencer.master_sequencer_D1046 =  pf_vf_mux_system_env_TB4_D1.master[146].sequencer;   
    sequencer.master_sequencer_D1047 =  pf_vf_mux_system_env_TB4_D1.master[147].sequencer;   
    sequencer.master_sequencer_D1048 =  pf_vf_mux_system_env_TB4_D1.master[148].sequencer;   
    sequencer.master_sequencer_D1049 =  pf_vf_mux_system_env_TB4_D1.master[149].sequencer;   
    sequencer.master_sequencer_D1050 =  pf_vf_mux_system_env_TB4_D1.master[150].sequencer;   
    sequencer.master_sequencer_D1051 =  pf_vf_mux_system_env_TB4_D1.master[151].sequencer;   
    sequencer.master_sequencer_D1052 =  pf_vf_mux_system_env_TB4_D1.master[152].sequencer;   
    sequencer.master_sequencer_D1053 =  pf_vf_mux_system_env_TB4_D1.master[153].sequencer;   
    sequencer.master_sequencer_D1054 =  pf_vf_mux_system_env_TB4_D1.master[154].sequencer;   
    sequencer.master_sequencer_D1055 =  pf_vf_mux_system_env_TB4_D1.master[155].sequencer;   
    sequencer.master_sequencer_D1056 =  pf_vf_mux_system_env_TB4_D1.master[156].sequencer;   
    sequencer.master_sequencer_D1057 =  pf_vf_mux_system_env_TB4_D1.master[157].sequencer;   
    sequencer.master_sequencer_D1058 =  pf_vf_mux_system_env_TB4_D1.master[158].sequencer;   
    sequencer.master_sequencer_D1059 =  pf_vf_mux_system_env_TB4_D1.master[159].sequencer;   
    sequencer.master_sequencer_D1060 =  pf_vf_mux_system_env_TB4_D1.master[160].sequencer;   
    sequencer.master_sequencer_D1061 =  pf_vf_mux_system_env_TB4_D1.master[161].sequencer;   
    sequencer.master_sequencer_D1062 =  pf_vf_mux_system_env_TB4_D1.master[162].sequencer;   
    sequencer.master_sequencer_D1063 =  pf_vf_mux_system_env_TB4_D1.master[163].sequencer;   
    sequencer.master_sequencer_D1064 =  pf_vf_mux_system_env_TB4_D1.master[164].sequencer;   
    sequencer.master_sequencer_D1065 =  pf_vf_mux_system_env_TB4_D1.master[165].sequencer;   
    sequencer.master_sequencer_D1066 =  pf_vf_mux_system_env_TB4_D1.master[166].sequencer;   
    sequencer.master_sequencer_D1067 =  pf_vf_mux_system_env_TB4_D1.master[167].sequencer;   
    sequencer.master_sequencer_D1068 =  pf_vf_mux_system_env_TB4_D1.master[168].sequencer;   
    sequencer.master_sequencer_D1069 =  pf_vf_mux_system_env_TB4_D1.master[169].sequencer;   
    sequencer.master_sequencer_D1070 =  pf_vf_mux_system_env_TB4_D1.master[170].sequencer;   
    sequencer.master_sequencer_D1071 =  pf_vf_mux_system_env_TB4_D1.master[171].sequencer;   
    sequencer.master_sequencer_D1072 =  pf_vf_mux_system_env_TB4_D1.master[172].sequencer;   
    sequencer.master_sequencer_D1073 =  pf_vf_mux_system_env_TB4_D1.master[173].sequencer;   
    sequencer.master_sequencer_D1074 =  pf_vf_mux_system_env_TB4_D1.master[174].sequencer;   
    sequencer.master_sequencer_D1075 =  pf_vf_mux_system_env_TB4_D1.master[175].sequencer;   
    sequencer.master_sequencer_D1076 =  pf_vf_mux_system_env_TB4_D1.master[176].sequencer;   
    sequencer.master_sequencer_D1077 =  pf_vf_mux_system_env_TB4_D1.master[177].sequencer;   
    sequencer.master_sequencer_D1078 =  pf_vf_mux_system_env_TB4_D1.master[178].sequencer;   
    sequencer.master_sequencer_D1079 =  pf_vf_mux_system_env_TB4_D1.master[179].sequencer;   
    sequencer.master_sequencer_D1080 =  pf_vf_mux_system_env_TB4_D1.master[180].sequencer;   
    sequencer.master_sequencer_D1081 =  pf_vf_mux_system_env_TB4_D1.master[181].sequencer;   
    sequencer.master_sequencer_D1082 =  pf_vf_mux_system_env_TB4_D1.master[182].sequencer;   
    sequencer.master_sequencer_D1083 =  pf_vf_mux_system_env_TB4_D1.master[183].sequencer;   
    sequencer.master_sequencer_D1084 =  pf_vf_mux_system_env_TB4_D1.master[184].sequencer;   
    sequencer.master_sequencer_D1085 =  pf_vf_mux_system_env_TB4_D1.master[185].sequencer;   
    sequencer.master_sequencer_D1086 =  pf_vf_mux_system_env_TB4_D1.master[186].sequencer;   
    sequencer.master_sequencer_D1087 =  pf_vf_mux_system_env_TB4_D1.master[187].sequencer;   
    sequencer.master_sequencer_D1088 =  pf_vf_mux_system_env_TB4_D1.master[188].sequencer;   
    sequencer.master_sequencer_D1089 =  pf_vf_mux_system_env_TB4_D1.master[189].sequencer;   
    sequencer.master_sequencer_D1090 =  pf_vf_mux_system_env_TB4_D1.master[190].sequencer;   
    sequencer.master_sequencer_D1091 =  pf_vf_mux_system_env_TB4_D1.master[191].sequencer;   
    sequencer.master_sequencer_D1092 =  pf_vf_mux_system_env_TB4_D1.master[192].sequencer;   
    sequencer.master_sequencer_D1093 =  pf_vf_mux_system_env_TB4_D1.master[193].sequencer;   
    sequencer.master_sequencer_D1094 =  pf_vf_mux_system_env_TB4_D1.master[194].sequencer;   
    sequencer.master_sequencer_D1095 =  pf_vf_mux_system_env_TB4_D1.master[195].sequencer;   
    sequencer.master_sequencer_D1096 =  pf_vf_mux_system_env_TB4_D1.master[196].sequencer;   
    sequencer.master_sequencer_D1097 =  pf_vf_mux_system_env_TB4_D1.master[197].sequencer;   
    sequencer.master_sequencer_D1098 =  pf_vf_mux_system_env_TB4_D1.master[198].sequencer;   
    sequencer.master_sequencer_D1099 =  pf_vf_mux_system_env_TB4_D1.master[199].sequencer;   
    sequencer.master_sequencer_D1100 =  pf_vf_mux_system_env_TB4_D1.master[200].sequencer;   
    sequencer.master_sequencer_D1101 =  pf_vf_mux_system_env_TB4_D1.master[201].sequencer;   
    sequencer.master_sequencer_D1102 =  pf_vf_mux_system_env_TB4_D1.master[202].sequencer;   
    sequencer.master_sequencer_D1103 =  pf_vf_mux_system_env_TB4_D1.master[203].sequencer;   
    sequencer.master_sequencer_D1104 =  pf_vf_mux_system_env_TB4_D1.master[204].sequencer;   
    sequencer.master_sequencer_D1105 =  pf_vf_mux_system_env_TB4_D1.master[205].sequencer;   
    sequencer.master_sequencer_D1106 =  pf_vf_mux_system_env_TB4_D1.master[206].sequencer;   
    sequencer.master_sequencer_D1107 =  pf_vf_mux_system_env_TB4_D1.master[207].sequencer;   
    sequencer.master_sequencer_D1108 =  pf_vf_mux_system_env_TB4_D1.master[208].sequencer;   
    sequencer.master_sequencer_D1109 =  pf_vf_mux_system_env_TB4_D1.master[209].sequencer;   
    sequencer.master_sequencer_D1110 =  pf_vf_mux_system_env_TB4_D1.master[210].sequencer;   
    sequencer.master_sequencer_D1111 =  pf_vf_mux_system_env_TB4_D1.master[211].sequencer;   
    sequencer.master_sequencer_D1112 =  pf_vf_mux_system_env_TB4_D1.master[212].sequencer;   
    sequencer.master_sequencer_D1113 =  pf_vf_mux_system_env_TB4_D1.master[213].sequencer;   
    sequencer.master_sequencer_D1114 =  pf_vf_mux_system_env_TB4_D1.master[214].sequencer;   
    sequencer.master_sequencer_D1115 =  pf_vf_mux_system_env_TB4_D1.master[215].sequencer;   
    sequencer.master_sequencer_D1116 =  pf_vf_mux_system_env_TB4_D1.master[216].sequencer;   
    sequencer.master_sequencer_D1117 =  pf_vf_mux_system_env_TB4_D1.master[217].sequencer;   
    sequencer.master_sequencer_D1118 =  pf_vf_mux_system_env_TB4_D1.master[218].sequencer;   
    sequencer.master_sequencer_D1119 =  pf_vf_mux_system_env_TB4_D1.master[219].sequencer;   
    sequencer.master_sequencer_D1120 =  pf_vf_mux_system_env_TB4_D1.master[220].sequencer;   
    sequencer.master_sequencer_D1121 =  pf_vf_mux_system_env_TB4_D1.master[221].sequencer;   
    sequencer.master_sequencer_D1122 =  pf_vf_mux_system_env_TB4_D1.master[222].sequencer;   
    sequencer.master_sequencer_D1123 =  pf_vf_mux_system_env_TB4_D1.master[223].sequencer;   
    sequencer.master_sequencer_D1124 =  pf_vf_mux_system_env_TB4_D1.master[224].sequencer;   
    sequencer.master_sequencer_D1125 =  pf_vf_mux_system_env_TB4_D1.master[225].sequencer;   
    sequencer.master_sequencer_D1126 =  pf_vf_mux_system_env_TB4_D1.master[226].sequencer;   
    sequencer.master_sequencer_D1127 =  pf_vf_mux_system_env_TB4_D1.master[227].sequencer;   
    sequencer.master_sequencer_D1128 =  pf_vf_mux_system_env_TB4_D1.master[228].sequencer;   
    sequencer.master_sequencer_D1129 =  pf_vf_mux_system_env_TB4_D1.master[229].sequencer;   
    sequencer.master_sequencer_D1130 =  pf_vf_mux_system_env_TB4_D1.master[230].sequencer;   
    sequencer.master_sequencer_D1131 =  pf_vf_mux_system_env_TB4_D1.master[231].sequencer;   
    sequencer.master_sequencer_D1132 =  pf_vf_mux_system_env_TB4_D1.master[232].sequencer;   
    sequencer.master_sequencer_D1133 =  pf_vf_mux_system_env_TB4_D1.master[233].sequencer;   
    sequencer.master_sequencer_D1134 =  pf_vf_mux_system_env_TB4_D1.master[234].sequencer;   
    sequencer.master_sequencer_D1135 =  pf_vf_mux_system_env_TB4_D1.master[235].sequencer;   
    sequencer.master_sequencer_D1136 =  pf_vf_mux_system_env_TB4_D1.master[236].sequencer;   
    sequencer.master_sequencer_D1137 =  pf_vf_mux_system_env_TB4_D1.master[237].sequencer;   
    sequencer.master_sequencer_D1138 =  pf_vf_mux_system_env_TB4_D1.master[238].sequencer;   
    sequencer.master_sequencer_D1139 =  pf_vf_mux_system_env_TB4_D1.master[239].sequencer;   
    sequencer.master_sequencer_D1140 =  pf_vf_mux_system_env_TB4_D1.master[240].sequencer;   
    sequencer.master_sequencer_D1141 =  pf_vf_mux_system_env_TB4_D1.master[241].sequencer;   
    sequencer.master_sequencer_D1142 =  pf_vf_mux_system_env_TB4_D1.master[242].sequencer;   
    sequencer.master_sequencer_D1143 =  pf_vf_mux_system_env_TB4_D1.master[243].sequencer;   
    sequencer.master_sequencer_D1144 =  pf_vf_mux_system_env_TB4_D1.master[244].sequencer;   
    sequencer.master_sequencer_D1145 =  pf_vf_mux_system_env_TB4_D1.master[245].sequencer;   
    sequencer.master_sequencer_D1146 =  pf_vf_mux_system_env_TB4_D1.master[246].sequencer;   
    sequencer.master_sequencer_D1147 =  pf_vf_mux_system_env_TB4_D1.master[247].sequencer;   
    sequencer.master_sequencer_D1148 =  pf_vf_mux_system_env_TB4_D1.master[248].sequencer;   
    sequencer.master_sequencer_D1149 =  pf_vf_mux_system_env_TB4_D1.master[249].sequencer;   
    sequencer.master_sequencer_D1150 =  pf_vf_mux_system_env_TB4_D1.master[250].sequencer;   
    sequencer.master_sequencer_D1151 =  pf_vf_mux_system_env_TB4_D1.master[251].sequencer;   
    sequencer.master_sequencer_D1152 =  pf_vf_mux_system_env_TB4_D1.master[252].sequencer;   
    sequencer.master_sequencer_D1153 =  pf_vf_mux_system_env_TB4_D1.master[253].sequencer;   
    sequencer.master_sequencer_D1154 =  pf_vf_mux_system_env_TB4_D1.master[254].sequencer;   
    sequencer.master_sequencer_D1155 =  pf_vf_mux_system_env_TB4_D1.master[255].sequencer;   
    sequencer.master_sequencer_D1156 =  pf_vf_mux_system_env_TB4_D1.master[256].sequencer;   
    sequencer.master_sequencer_D1157 =  pf_vf_mux_system_env_TB4_D1.master[257].sequencer;   
    sequencer.master_sequencer_D1158 =  pf_vf_mux_system_env_TB4_D1.master[258].sequencer;   
    sequencer.master_sequencer_D1159 =  pf_vf_mux_system_env_TB4_D1.master[259].sequencer;   
    sequencer.master_sequencer_D1160 =  pf_vf_mux_system_env_TB4_D1.master[260].sequencer;   
    sequencer.master_sequencer_D1161 =  pf_vf_mux_system_env_TB4_D1.master[261].sequencer;   
    sequencer.master_sequencer_D1162 =  pf_vf_mux_system_env_TB4_D1.master[262].sequencer;   
    sequencer.master_sequencer_D1163 =  pf_vf_mux_system_env_TB4_D1.master[263].sequencer;   
    sequencer.master_sequencer_D1164 =  pf_vf_mux_system_env_TB4_D1.master[264].sequencer;   
    sequencer.master_sequencer_D1165 =  pf_vf_mux_system_env_TB4_D1.master[265].sequencer;   
    sequencer.master_sequencer_D1166 =  pf_vf_mux_system_env_TB4_D1.master[266].sequencer;   
    sequencer.master_sequencer_D1167 =  pf_vf_mux_system_env_TB4_D1.master[267].sequencer;   
    sequencer.master_sequencer_D1168 =  pf_vf_mux_system_env_TB4_D1.master[268].sequencer;   
    sequencer.master_sequencer_D1169 =  pf_vf_mux_system_env_TB4_D1.master[269].sequencer;   
    sequencer.master_sequencer_D1170 =  pf_vf_mux_system_env_TB4_D1.master[270].sequencer;   
    sequencer.master_sequencer_D1171 =  pf_vf_mux_system_env_TB4_D1.master[271].sequencer;   
    sequencer.master_sequencer_D1172 =  pf_vf_mux_system_env_TB4_D1.master[272].sequencer;   
    sequencer.master_sequencer_D1173 =  pf_vf_mux_system_env_TB4_D1.master[273].sequencer;   
    sequencer.master_sequencer_D1174 =  pf_vf_mux_system_env_TB4_D1.master[274].sequencer;   
    sequencer.master_sequencer_D1175 =  pf_vf_mux_system_env_TB4_D1.master[275].sequencer;   
    sequencer.master_sequencer_D1176 =  pf_vf_mux_system_env_TB4_D1.master[276].sequencer;   
    sequencer.master_sequencer_D1177 =  pf_vf_mux_system_env_TB4_D1.master[277].sequencer;   
    sequencer.master_sequencer_D1178 =  pf_vf_mux_system_env_TB4_D1.master[278].sequencer;   
    sequencer.master_sequencer_D1179 =  pf_vf_mux_system_env_TB4_D1.master[279].sequencer;   
    sequencer.master_sequencer_D1180 =  pf_vf_mux_system_env_TB4_D1.master[280].sequencer;   
    sequencer.master_sequencer_D1181 =  pf_vf_mux_system_env_TB4_D1.master[281].sequencer;   
    sequencer.master_sequencer_D1182 =  pf_vf_mux_system_env_TB4_D1.master[282].sequencer;   
    sequencer.master_sequencer_D1183 =  pf_vf_mux_system_env_TB4_D1.master[283].sequencer;   
    sequencer.master_sequencer_D1184 =  pf_vf_mux_system_env_TB4_D1.master[284].sequencer;   
    sequencer.master_sequencer_D1185 =  pf_vf_mux_system_env_TB4_D1.master[285].sequencer;   
    sequencer.master_sequencer_D1186 =  pf_vf_mux_system_env_TB4_D1.master[286].sequencer;   
    sequencer.master_sequencer_D1187 =  pf_vf_mux_system_env_TB4_D1.master[287].sequencer;   
    sequencer.master_sequencer_D1188 =  pf_vf_mux_system_env_TB4_D1.master[288].sequencer;   
    sequencer.master_sequencer_D1189 =  pf_vf_mux_system_env_TB4_D1.master[289].sequencer;   
    sequencer.master_sequencer_D1190 =  pf_vf_mux_system_env_TB4_D1.master[290].sequencer;   
    sequencer.master_sequencer_D1191 =  pf_vf_mux_system_env_TB4_D1.master[291].sequencer;   
    sequencer.master_sequencer_D1192 =  pf_vf_mux_system_env_TB4_D1.master[292].sequencer;   
    sequencer.master_sequencer_D1193 =  pf_vf_mux_system_env_TB4_D1.master[293].sequencer;   
    sequencer.master_sequencer_D1194 =  pf_vf_mux_system_env_TB4_D1.master[294].sequencer;   
    sequencer.master_sequencer_D1195 =  pf_vf_mux_system_env_TB4_D1.master[295].sequencer;   
    sequencer.master_sequencer_D1196 =  pf_vf_mux_system_env_TB4_D1.master[296].sequencer;   
    sequencer.master_sequencer_D1197 =  pf_vf_mux_system_env_TB4_D1.master[297].sequencer;   
    sequencer.master_sequencer_D1198 =  pf_vf_mux_system_env_TB4_D1.master[298].sequencer;   
    sequencer.master_sequencer_D1199 =  pf_vf_mux_system_env_TB4_D1.master[299].sequencer;   
    sequencer.master_sequencer_D1200 =  pf_vf_mux_system_env_TB4_D1.master[300].sequencer;   
    sequencer.master_sequencer_D1201 =  pf_vf_mux_system_env_TB4_D1.master[301].sequencer;   
    sequencer.master_sequencer_D1202 =  pf_vf_mux_system_env_TB4_D1.master[302].sequencer;   
    sequencer.master_sequencer_D1203 =  pf_vf_mux_system_env_TB4_D1.master[303].sequencer;   
    sequencer.master_sequencer_D1204 =  pf_vf_mux_system_env_TB4_D1.master[304].sequencer;   
    sequencer.master_sequencer_D1205 =  pf_vf_mux_system_env_TB4_D1.master[305].sequencer;   
    sequencer.master_sequencer_D1206 =  pf_vf_mux_system_env_TB4_D1.master[306].sequencer;   
    sequencer.master_sequencer_D1207 =  pf_vf_mux_system_env_TB4_D1.master[307].sequencer;   
    sequencer.master_sequencer_D1208 =  pf_vf_mux_system_env_TB4_D1.master[308].sequencer;   
    sequencer.master_sequencer_D1209 =  pf_vf_mux_system_env_TB4_D1.master[309].sequencer;   
    sequencer.master_sequencer_D1210 =  pf_vf_mux_system_env_TB4_D1.master[310].sequencer;   
    sequencer.master_sequencer_D1211 =  pf_vf_mux_system_env_TB4_D1.master[311].sequencer;   
    sequencer.master_sequencer_D1212 =  pf_vf_mux_system_env_TB4_D1.master[312].sequencer;   
    sequencer.master_sequencer_D1213 =  pf_vf_mux_system_env_TB4_D1.master[313].sequencer;   
    sequencer.master_sequencer_D1214 =  pf_vf_mux_system_env_TB4_D1.master[314].sequencer;   
    sequencer.master_sequencer_D1215 =  pf_vf_mux_system_env_TB4_D1.master[315].sequencer;   
    sequencer.master_sequencer_D1216 =  pf_vf_mux_system_env_TB4_D1.master[316].sequencer;   
    sequencer.master_sequencer_D1217 =  pf_vf_mux_system_env_TB4_D1.master[317].sequencer;   
    sequencer.master_sequencer_D1218 =  pf_vf_mux_system_env_TB4_D1.master[318].sequencer;   
    sequencer.master_sequencer_D1219 =  pf_vf_mux_system_env_TB4_D1.master[319].sequencer;   
    sequencer.master_sequencer_D1220 =  pf_vf_mux_system_env_TB4_D1.master[320].sequencer;   
    sequencer.master_sequencer_D1221 =  pf_vf_mux_system_env_TB4_D1.master[321].sequencer;   
    sequencer.master_sequencer_D1222 =  pf_vf_mux_system_env_TB4_D1.master[322].sequencer;   
    sequencer.master_sequencer_D1223 =  pf_vf_mux_system_env_TB4_D1.master[323].sequencer;   
    sequencer.master_sequencer_D1224 =  pf_vf_mux_system_env_TB4_D1.master[324].sequencer;   
    sequencer.master_sequencer_D1225 =  pf_vf_mux_system_env_TB4_D1.master[325].sequencer;   
    sequencer.master_sequencer_D1226 =  pf_vf_mux_system_env_TB4_D1.master[326].sequencer;   
    sequencer.master_sequencer_D1227 =  pf_vf_mux_system_env_TB4_D1.master[327].sequencer;   
    sequencer.master_sequencer_D1228 =  pf_vf_mux_system_env_TB4_D1.master[328].sequencer;   
    sequencer.master_sequencer_D1229 =  pf_vf_mux_system_env_TB4_D1.master[329].sequencer;   
    sequencer.master_sequencer_D1230 =  pf_vf_mux_system_env_TB4_D1.master[330].sequencer;   
    sequencer.master_sequencer_D1231 =  pf_vf_mux_system_env_TB4_D1.master[331].sequencer;   
    sequencer.master_sequencer_D1232 =  pf_vf_mux_system_env_TB4_D1.master[332].sequencer;   
    sequencer.master_sequencer_D1233 =  pf_vf_mux_system_env_TB4_D1.master[333].sequencer;   
    sequencer.master_sequencer_D1234 =  pf_vf_mux_system_env_TB4_D1.master[334].sequencer;   
    sequencer.master_sequencer_D1235 =  pf_vf_mux_system_env_TB4_D1.master[335].sequencer;   
    sequencer.master_sequencer_D1236 =  pf_vf_mux_system_env_TB4_D1.master[336].sequencer;   
    sequencer.master_sequencer_D1237 =  pf_vf_mux_system_env_TB4_D1.master[337].sequencer;   
    sequencer.master_sequencer_D1238 =  pf_vf_mux_system_env_TB4_D1.master[338].sequencer;   
    sequencer.master_sequencer_D1239 =  pf_vf_mux_system_env_TB4_D1.master[339].sequencer;   
    sequencer.master_sequencer_D1240 =  pf_vf_mux_system_env_TB4_D1.master[340].sequencer;   
    sequencer.master_sequencer_D1241 =  pf_vf_mux_system_env_TB4_D1.master[341].sequencer;   
    sequencer.master_sequencer_D1242 =  pf_vf_mux_system_env_TB4_D1.master[342].sequencer;   
    sequencer.master_sequencer_D1243 =  pf_vf_mux_system_env_TB4_D1.master[343].sequencer;   
    sequencer.master_sequencer_D1244 =  pf_vf_mux_system_env_TB4_D1.master[344].sequencer;   
    sequencer.master_sequencer_D1245 =  pf_vf_mux_system_env_TB4_D1.master[345].sequencer;   
    sequencer.master_sequencer_D1246 =  pf_vf_mux_system_env_TB4_D1.master[346].sequencer;   
    sequencer.master_sequencer_D1247 =  pf_vf_mux_system_env_TB4_D1.master[347].sequencer;   
    sequencer.master_sequencer_D1248 =  pf_vf_mux_system_env_TB4_D1.master[348].sequencer;   
    sequencer.master_sequencer_D1249 =  pf_vf_mux_system_env_TB4_D1.master[349].sequencer;   
    sequencer.master_sequencer_D1250 =  pf_vf_mux_system_env_TB4_D1.master[350].sequencer;   
    sequencer.master_sequencer_D1251 =  pf_vf_mux_system_env_TB4_D1.master[351].sequencer;   
    sequencer.master_sequencer_D1252 =  pf_vf_mux_system_env_TB4_D1.master[352].sequencer;   
    sequencer.master_sequencer_D1253 =  pf_vf_mux_system_env_TB4_D1.master[353].sequencer;   
    sequencer.master_sequencer_D1254 =  pf_vf_mux_system_env_TB4_D1.master[354].sequencer;   
    sequencer.master_sequencer_D1255 =  pf_vf_mux_system_env_TB4_D1.master[355].sequencer;   
    sequencer.master_sequencer_D1256 =  pf_vf_mux_system_env_TB4_D1.master[356].sequencer;   
    sequencer.master_sequencer_D1257 =  pf_vf_mux_system_env_TB4_D1.master[357].sequencer;   
    sequencer.master_sequencer_D1258 =  pf_vf_mux_system_env_TB4_D1.master[358].sequencer;   
    sequencer.master_sequencer_D1259 =  pf_vf_mux_system_env_TB4_D1.master[359].sequencer;   
    sequencer.master_sequencer_D1260 =  pf_vf_mux_system_env_TB4_D1.master[360].sequencer;   
    sequencer.master_sequencer_D1261 =  pf_vf_mux_system_env_TB4_D1.master[361].sequencer;   
    sequencer.master_sequencer_D1262 =  pf_vf_mux_system_env_TB4_D1.master[362].sequencer;   
    sequencer.master_sequencer_D1263 =  pf_vf_mux_system_env_TB4_D1.master[363].sequencer;   
    sequencer.master_sequencer_D1264 =  pf_vf_mux_system_env_TB4_D1.master[364].sequencer;   
    sequencer.master_sequencer_D1265 =  pf_vf_mux_system_env_TB4_D1.master[365].sequencer;   
    sequencer.master_sequencer_D1266 =  pf_vf_mux_system_env_TB4_D1.master[366].sequencer;   
    sequencer.master_sequencer_D1267 =  pf_vf_mux_system_env_TB4_D1.master[367].sequencer;   
    sequencer.master_sequencer_D1268 =  pf_vf_mux_system_env_TB4_D1.master[368].sequencer;   
    sequencer.master_sequencer_D1269 =  pf_vf_mux_system_env_TB4_D1.master[369].sequencer;   
    sequencer.master_sequencer_D1270 =  pf_vf_mux_system_env_TB4_D1.master[370].sequencer;   
    sequencer.master_sequencer_D1271 =  pf_vf_mux_system_env_TB4_D1.master[371].sequencer;   
    sequencer.master_sequencer_D1272 =  pf_vf_mux_system_env_TB4_D1.master[372].sequencer;   
    sequencer.master_sequencer_D1273 =  pf_vf_mux_system_env_TB4_D1.master[373].sequencer;   
    sequencer.master_sequencer_D1274 =  pf_vf_mux_system_env_TB4_D1.master[374].sequencer;   
    sequencer.master_sequencer_D1275 =  pf_vf_mux_system_env_TB4_D1.master[375].sequencer;   
    sequencer.master_sequencer_D1276 =  pf_vf_mux_system_env_TB4_D1.master[376].sequencer;   
    sequencer.master_sequencer_D1277 =  pf_vf_mux_system_env_TB4_D1.master[377].sequencer;   
    sequencer.master_sequencer_D1278 =  pf_vf_mux_system_env_TB4_D1.master[378].sequencer;   
    sequencer.master_sequencer_D1279 =  pf_vf_mux_system_env_TB4_D1.master[379].sequencer;   
    sequencer.master_sequencer_D1280 =  pf_vf_mux_system_env_TB4_D1.master[380].sequencer;   
    sequencer.master_sequencer_D1281 =  pf_vf_mux_system_env_TB4_D1.master[381].sequencer;   
    sequencer.master_sequencer_D1282 =  pf_vf_mux_system_env_TB4_D1.master[382].sequencer;   
    sequencer.master_sequencer_D1283 =  pf_vf_mux_system_env_TB4_D1.master[383].sequencer;   
    sequencer.master_sequencer_D1284 =  pf_vf_mux_system_env_TB4_D1.master[384].sequencer;   
    sequencer.master_sequencer_D1285 =  pf_vf_mux_system_env_TB4_D1.master[385].sequencer;   
    sequencer.master_sequencer_D1286 =  pf_vf_mux_system_env_TB4_D1.master[386].sequencer;   
    sequencer.master_sequencer_D1287 =  pf_vf_mux_system_env_TB4_D1.master[387].sequencer;   
    sequencer.master_sequencer_D1288 =  pf_vf_mux_system_env_TB4_D1.master[388].sequencer;   
    sequencer.master_sequencer_D1289 =  pf_vf_mux_system_env_TB4_D1.master[389].sequencer;   
    sequencer.master_sequencer_D1290 =  pf_vf_mux_system_env_TB4_D1.master[390].sequencer;   
    sequencer.master_sequencer_D1291 =  pf_vf_mux_system_env_TB4_D1.master[391].sequencer;   
    sequencer.master_sequencer_D1292 =  pf_vf_mux_system_env_TB4_D1.master[392].sequencer;   
    sequencer.master_sequencer_D1293 =  pf_vf_mux_system_env_TB4_D1.master[393].sequencer;   
    sequencer.master_sequencer_D1294 =  pf_vf_mux_system_env_TB4_D1.master[394].sequencer;   
    sequencer.master_sequencer_D1295 =  pf_vf_mux_system_env_TB4_D1.master[395].sequencer;   
    sequencer.master_sequencer_D1296 =  pf_vf_mux_system_env_TB4_D1.master[396].sequencer;   
    sequencer.master_sequencer_D1297 =  pf_vf_mux_system_env_TB4_D1.master[397].sequencer;   
    sequencer.master_sequencer_D1298 =  pf_vf_mux_system_env_TB4_D1.master[398].sequencer;   
    sequencer.master_sequencer_D1299 =  pf_vf_mux_system_env_TB4_D1.master[399].sequencer;   
    sequencer.master_sequencer_D1300 =  pf_vf_mux_system_env_TB4_D1.master[400].sequencer;   
    sequencer.master_sequencer_D1301 =  pf_vf_mux_system_env_TB4_D1.master[401].sequencer;   
    sequencer.master_sequencer_D1302 =  pf_vf_mux_system_env_TB4_D1.master[402].sequencer;   
    sequencer.master_sequencer_D1303 =  pf_vf_mux_system_env_TB4_D1.master[403].sequencer;   
    sequencer.master_sequencer_D1304 =  pf_vf_mux_system_env_TB4_D1.master[404].sequencer;   
    sequencer.master_sequencer_D1305 =  pf_vf_mux_system_env_TB4_D1.master[405].sequencer;   
    sequencer.master_sequencer_D1306 =  pf_vf_mux_system_env_TB4_D1.master[406].sequencer;   
    sequencer.master_sequencer_D1307 =  pf_vf_mux_system_env_TB4_D1.master[407].sequencer;   
    sequencer.master_sequencer_D1308 =  pf_vf_mux_system_env_TB4_D1.master[408].sequencer;   
    sequencer.master_sequencer_D1309 =  pf_vf_mux_system_env_TB4_D1.master[409].sequencer;   
    sequencer.master_sequencer_D1310 =  pf_vf_mux_system_env_TB4_D1.master[410].sequencer;   
    sequencer.master_sequencer_D1311 =  pf_vf_mux_system_env_TB4_D1.master[411].sequencer;   
    sequencer.master_sequencer_D1312 =  pf_vf_mux_system_env_TB4_D1.master[412].sequencer;   
    sequencer.master_sequencer_D1313 =  pf_vf_mux_system_env_TB4_D1.master[413].sequencer;   
    sequencer.master_sequencer_D1314 =  pf_vf_mux_system_env_TB4_D1.master[414].sequencer;   
    sequencer.master_sequencer_D1315 =  pf_vf_mux_system_env_TB4_D1.master[415].sequencer;   
    sequencer.master_sequencer_D1316 =  pf_vf_mux_system_env_TB4_D1.master[416].sequencer;   
    sequencer.master_sequencer_D1317 =  pf_vf_mux_system_env_TB4_D1.master[417].sequencer;   
    sequencer.master_sequencer_D1318 =  pf_vf_mux_system_env_TB4_D1.master[418].sequencer;   
    sequencer.master_sequencer_D1319 =  pf_vf_mux_system_env_TB4_D1.master[419].sequencer;   
    sequencer.master_sequencer_D1320 =  pf_vf_mux_system_env_TB4_D1.master[420].sequencer;   
    sequencer.master_sequencer_D1321 =  pf_vf_mux_system_env_TB4_D1.master[421].sequencer;   
    sequencer.master_sequencer_D1322 =  pf_vf_mux_system_env_TB4_D1.master[422].sequencer;   
    sequencer.master_sequencer_D1323 =  pf_vf_mux_system_env_TB4_D1.master[423].sequencer;   
    sequencer.master_sequencer_D1324 =  pf_vf_mux_system_env_TB4_D1.master[424].sequencer;   
    sequencer.master_sequencer_D1325 =  pf_vf_mux_system_env_TB4_D1.master[425].sequencer;   
    sequencer.master_sequencer_D1326 =  pf_vf_mux_system_env_TB4_D1.master[426].sequencer;   
    sequencer.master_sequencer_D1327 =  pf_vf_mux_system_env_TB4_D1.master[427].sequencer;   
    sequencer.master_sequencer_D1328 =  pf_vf_mux_system_env_TB4_D1.master[428].sequencer;   
    sequencer.master_sequencer_D1329 =  pf_vf_mux_system_env_TB4_D1.master[429].sequencer;   
    sequencer.master_sequencer_D1330 =  pf_vf_mux_system_env_TB4_D1.master[430].sequencer;   
    sequencer.master_sequencer_D1331 =  pf_vf_mux_system_env_TB4_D1.master[431].sequencer;   
    sequencer.master_sequencer_D1332 =  pf_vf_mux_system_env_TB4_D1.master[432].sequencer;   
    sequencer.master_sequencer_D1333 =  pf_vf_mux_system_env_TB4_D1.master[433].sequencer;   
    sequencer.master_sequencer_D1334 =  pf_vf_mux_system_env_TB4_D1.master[434].sequencer;   
    sequencer.master_sequencer_D1335 =  pf_vf_mux_system_env_TB4_D1.master[435].sequencer;   
    sequencer.master_sequencer_D1336 =  pf_vf_mux_system_env_TB4_D1.master[436].sequencer;   
    sequencer.master_sequencer_D1337 =  pf_vf_mux_system_env_TB4_D1.master[437].sequencer;   
    sequencer.master_sequencer_D1338 =  pf_vf_mux_system_env_TB4_D1.master[438].sequencer;   
    sequencer.master_sequencer_D1339 =  pf_vf_mux_system_env_TB4_D1.master[439].sequencer;   
    sequencer.master_sequencer_D1340 =  pf_vf_mux_system_env_TB4_D1.master[440].sequencer;   
    sequencer.master_sequencer_D1341 =  pf_vf_mux_system_env_TB4_D1.master[441].sequencer;   
    sequencer.master_sequencer_D1342 =  pf_vf_mux_system_env_TB4_D1.master[442].sequencer;   
    sequencer.master_sequencer_D1343 =  pf_vf_mux_system_env_TB4_D1.master[443].sequencer;   
    sequencer.master_sequencer_D1344 =  pf_vf_mux_system_env_TB4_D1.master[444].sequencer;   
    sequencer.master_sequencer_D1345 =  pf_vf_mux_system_env_TB4_D1.master[445].sequencer;   
    sequencer.master_sequencer_D1346 =  pf_vf_mux_system_env_TB4_D1.master[446].sequencer;   
    sequencer.master_sequencer_D1347 =  pf_vf_mux_system_env_TB4_D1.master[447].sequencer;   
    sequencer.master_sequencer_D1348 =  pf_vf_mux_system_env_TB4_D1.master[448].sequencer;   
    sequencer.master_sequencer_D1349 =  pf_vf_mux_system_env_TB4_D1.master[449].sequencer;
    sequencer.master_sequencer_D1350 =  pf_vf_mux_system_env_TB4_D2.master[0].sequencer;   
    sequencer.master_sequencer_D1351 =  pf_vf_mux_system_env_TB4_D2.master[1].sequencer;   
    sequencer.master_sequencer_D1352 =  pf_vf_mux_system_env_TB4_D2.master[2].sequencer;   
    sequencer.master_sequencer_D1353 =  pf_vf_mux_system_env_TB4_D2.master[3].sequencer;   
    sequencer.master_sequencer_D1354 =  pf_vf_mux_system_env_TB4_D2.master[4].sequencer;   
    sequencer.master_sequencer_D1355 =  pf_vf_mux_system_env_TB4_D2.master[5].sequencer;   
    sequencer.master_sequencer_D1356 =  pf_vf_mux_system_env_TB4_D2.master[6].sequencer;   
    sequencer.master_sequencer_D1357 =  pf_vf_mux_system_env_TB4_D2.master[7].sequencer;   
    sequencer.master_sequencer_D1358 =  pf_vf_mux_system_env_TB4_D2.master[8].sequencer;   
    sequencer.master_sequencer_D1359 =  pf_vf_mux_system_env_TB4_D2.master[9].sequencer;   
    sequencer.master_sequencer_D1360 =  pf_vf_mux_system_env_TB4_D2.master[10].sequencer;   
    sequencer.master_sequencer_D1361 =  pf_vf_mux_system_env_TB4_D2.master[11].sequencer;   
    sequencer.master_sequencer_D1362 =  pf_vf_mux_system_env_TB4_D2.master[12].sequencer;   
    sequencer.master_sequencer_D1363 =  pf_vf_mux_system_env_TB4_D2.master[13].sequencer;   
    sequencer.master_sequencer_D1364 =  pf_vf_mux_system_env_TB4_D2.master[14].sequencer;   
    sequencer.master_sequencer_D1365 =  pf_vf_mux_system_env_TB4_D2.master[15].sequencer;   
    sequencer.master_sequencer_D1366 =  pf_vf_mux_system_env_TB4_D2.master[16].sequencer;   
    sequencer.master_sequencer_D1367 =  pf_vf_mux_system_env_TB4_D2.master[17].sequencer;   
    sequencer.master_sequencer_D1368 =  pf_vf_mux_system_env_TB4_D2.master[18].sequencer;   
    sequencer.master_sequencer_D1369 =  pf_vf_mux_system_env_TB4_D2.master[19].sequencer;   
    sequencer.master_sequencer_D1370 =  pf_vf_mux_system_env_TB4_D2.master[20].sequencer;   
    sequencer.master_sequencer_D1371 =  pf_vf_mux_system_env_TB4_D2.master[21].sequencer;   
    sequencer.master_sequencer_D1372 =  pf_vf_mux_system_env_TB4_D2.master[22].sequencer;   
    sequencer.master_sequencer_D1373 =  pf_vf_mux_system_env_TB4_D2.master[23].sequencer;   
    sequencer.master_sequencer_D1374 =  pf_vf_mux_system_env_TB4_D2.master[24].sequencer;   
    sequencer.master_sequencer_D1375 =  pf_vf_mux_system_env_TB4_D2.master[25].sequencer;   
    sequencer.master_sequencer_D1376 =  pf_vf_mux_system_env_TB4_D2.master[26].sequencer;   
    sequencer.master_sequencer_D1377 =  pf_vf_mux_system_env_TB4_D2.master[27].sequencer;   
    sequencer.master_sequencer_D1378 =  pf_vf_mux_system_env_TB4_D2.master[28].sequencer;   
    sequencer.master_sequencer_D1379 =  pf_vf_mux_system_env_TB4_D2.master[29].sequencer;   
    sequencer.master_sequencer_D1380 =  pf_vf_mux_system_env_TB4_D2.master[30].sequencer;   
    sequencer.master_sequencer_D1381 =  pf_vf_mux_system_env_TB4_D2.master[31].sequencer;   
    sequencer.master_sequencer_D1382 =  pf_vf_mux_system_env_TB4_D2.master[32].sequencer;   
    sequencer.master_sequencer_D1383 =  pf_vf_mux_system_env_TB4_D2.master[33].sequencer;   
    sequencer.master_sequencer_D1384 =  pf_vf_mux_system_env_TB4_D2.master[34].sequencer;   
    sequencer.master_sequencer_D1385 =  pf_vf_mux_system_env_TB4_D2.master[35].sequencer;   
    sequencer.master_sequencer_D1386 =  pf_vf_mux_system_env_TB4_D2.master[36].sequencer;   
    sequencer.master_sequencer_D1387 =  pf_vf_mux_system_env_TB4_D2.master[37].sequencer;   
    sequencer.master_sequencer_D1388 =  pf_vf_mux_system_env_TB4_D2.master[38].sequencer;   
    sequencer.master_sequencer_D1389 =  pf_vf_mux_system_env_TB4_D2.master[39].sequencer;   
    sequencer.master_sequencer_D1390 =  pf_vf_mux_system_env_TB4_D2.master[40].sequencer;   
    sequencer.master_sequencer_D1391 =  pf_vf_mux_system_env_TB4_D2.master[41].sequencer;   
    sequencer.master_sequencer_D1392 =  pf_vf_mux_system_env_TB4_D2.master[42].sequencer;   
    sequencer.master_sequencer_D1393 =  pf_vf_mux_system_env_TB4_D2.master[43].sequencer;   
    sequencer.master_sequencer_D1394 =  pf_vf_mux_system_env_TB4_D2.master[44].sequencer;   
    sequencer.master_sequencer_D1395 =  pf_vf_mux_system_env_TB4_D2.master[45].sequencer;   
    sequencer.master_sequencer_D1396 =  pf_vf_mux_system_env_TB4_D2.master[46].sequencer;   
    sequencer.master_sequencer_D1397 =  pf_vf_mux_system_env_TB4_D2.master[47].sequencer;   
    sequencer.master_sequencer_D1398 =  pf_vf_mux_system_env_TB4_D2.master[48].sequencer;   
    sequencer.master_sequencer_D1399 =  pf_vf_mux_system_env_TB4_D2.master[49].sequencer;   
    sequencer.master_sequencer_D1400 =  pf_vf_mux_system_env_TB4_D2.master[50].sequencer;   
    sequencer.master_sequencer_D1401 =  pf_vf_mux_system_env_TB4_D2.master[51].sequencer;   
    sequencer.master_sequencer_D1402 =  pf_vf_mux_system_env_TB4_D2.master[52].sequencer;   
    sequencer.master_sequencer_D1403 =  pf_vf_mux_system_env_TB4_D2.master[53].sequencer;   
    sequencer.master_sequencer_D1404 =  pf_vf_mux_system_env_TB4_D2.master[54].sequencer;   
    sequencer.master_sequencer_D1405 =  pf_vf_mux_system_env_TB4_D2.master[55].sequencer;   
    sequencer.master_sequencer_D1406 =  pf_vf_mux_system_env_TB4_D2.master[56].sequencer;   
    sequencer.master_sequencer_D1407 =  pf_vf_mux_system_env_TB4_D2.master[57].sequencer;   
    sequencer.master_sequencer_D1408 =  pf_vf_mux_system_env_TB4_D2.master[58].sequencer;   
    sequencer.master_sequencer_D1409 =  pf_vf_mux_system_env_TB4_D2.master[59].sequencer;   
    sequencer.master_sequencer_D1410 =  pf_vf_mux_system_env_TB4_D2.master[60].sequencer;   
    sequencer.master_sequencer_D1411 =  pf_vf_mux_system_env_TB4_D2.master[61].sequencer;   
    sequencer.master_sequencer_D1412 =  pf_vf_mux_system_env_TB4_D2.master[62].sequencer;   
    sequencer.master_sequencer_D1413 =  pf_vf_mux_system_env_TB4_D2.master[63].sequencer;   
    sequencer.master_sequencer_D1414 =  pf_vf_mux_system_env_TB4_D2.master[64].sequencer;   
    sequencer.master_sequencer_D1415 =  pf_vf_mux_system_env_TB4_D2.master[65].sequencer;   
    sequencer.master_sequencer_D1416 =  pf_vf_mux_system_env_TB4_D2.master[66].sequencer;   
    sequencer.master_sequencer_D1417 =  pf_vf_mux_system_env_TB4_D2.master[67].sequencer;   
    sequencer.master_sequencer_D1418 =  pf_vf_mux_system_env_TB4_D2.master[68].sequencer;   
    sequencer.master_sequencer_D1419 =  pf_vf_mux_system_env_TB4_D2.master[69].sequencer;   
    sequencer.master_sequencer_D1420 =  pf_vf_mux_system_env_TB4_D2.master[70].sequencer;   
    sequencer.master_sequencer_D1421 =  pf_vf_mux_system_env_TB4_D2.master[71].sequencer;   
    sequencer.master_sequencer_D1422 =  pf_vf_mux_system_env_TB4_D2.master[72].sequencer;   
    sequencer.master_sequencer_D1423 =  pf_vf_mux_system_env_TB4_D2.master[73].sequencer;   
    sequencer.master_sequencer_D1424 =  pf_vf_mux_system_env_TB4_D2.master[74].sequencer;   
    sequencer.master_sequencer_D1425 =  pf_vf_mux_system_env_TB4_D2.master[75].sequencer;   
    sequencer.master_sequencer_D1426 =  pf_vf_mux_system_env_TB4_D2.master[76].sequencer;   
    sequencer.master_sequencer_D1427 =  pf_vf_mux_system_env_TB4_D2.master[77].sequencer;   
    sequencer.master_sequencer_D1428 =  pf_vf_mux_system_env_TB4_D2.master[78].sequencer;   
    sequencer.master_sequencer_D1429 =  pf_vf_mux_system_env_TB4_D2.master[79].sequencer;   
    sequencer.master_sequencer_D1430 =  pf_vf_mux_system_env_TB4_D2.master[80].sequencer;   
    sequencer.master_sequencer_D1431 =  pf_vf_mux_system_env_TB4_D2.master[81].sequencer;   
    sequencer.master_sequencer_D1432 =  pf_vf_mux_system_env_TB4_D2.master[82].sequencer;   
    sequencer.master_sequencer_D1433 =  pf_vf_mux_system_env_TB4_D2.master[83].sequencer;   
    sequencer.master_sequencer_D1434 =  pf_vf_mux_system_env_TB4_D2.master[84].sequencer;   
    sequencer.master_sequencer_D1435 =  pf_vf_mux_system_env_TB4_D2.master[85].sequencer;   
    sequencer.master_sequencer_D1436 =  pf_vf_mux_system_env_TB4_D2.master[86].sequencer;   
    sequencer.master_sequencer_D1437 =  pf_vf_mux_system_env_TB4_D2.master[87].sequencer;   
    sequencer.master_sequencer_D1438 =  pf_vf_mux_system_env_TB4_D2.master[88].sequencer;   
    sequencer.master_sequencer_D1439 =  pf_vf_mux_system_env_TB4_D2.master[89].sequencer;   
    sequencer.master_sequencer_D1440 =  pf_vf_mux_system_env_TB4_D2.master[90].sequencer;   
    sequencer.master_sequencer_D1441 =  pf_vf_mux_system_env_TB4_D2.master[91].sequencer;   
    sequencer.master_sequencer_D1442 =  pf_vf_mux_system_env_TB4_D2.master[92].sequencer;   
    sequencer.master_sequencer_D1443 =  pf_vf_mux_system_env_TB4_D2.master[93].sequencer;   
    sequencer.master_sequencer_D1444 =  pf_vf_mux_system_env_TB4_D2.master[94].sequencer;   
    sequencer.master_sequencer_D1445 =  pf_vf_mux_system_env_TB4_D2.master[95].sequencer;   
    sequencer.master_sequencer_D1446 =  pf_vf_mux_system_env_TB4_D2.master[96].sequencer;   
    sequencer.master_sequencer_D1447 =  pf_vf_mux_system_env_TB4_D2.master[97].sequencer;   
    sequencer.master_sequencer_D1448 =  pf_vf_mux_system_env_TB4_D2.master[98].sequencer;   
    sequencer.master_sequencer_D1449 =  pf_vf_mux_system_env_TB4_D2.master[99].sequencer;   
    sequencer.master_sequencer_D1450 =  pf_vf_mux_system_env_TB4_D2.master[100].sequencer;   
    sequencer.master_sequencer_D1451 =  pf_vf_mux_system_env_TB4_D2.master[101].sequencer;   
    sequencer.master_sequencer_D1452 =  pf_vf_mux_system_env_TB4_D2.master[102].sequencer;   
    sequencer.master_sequencer_D1453 =  pf_vf_mux_system_env_TB4_D2.master[103].sequencer;   
    sequencer.master_sequencer_D1454 =  pf_vf_mux_system_env_TB4_D2.master[104].sequencer;   
    sequencer.master_sequencer_D1455 =  pf_vf_mux_system_env_TB4_D2.master[105].sequencer;   
    sequencer.master_sequencer_D1456 =  pf_vf_mux_system_env_TB4_D2.master[106].sequencer;   
    sequencer.master_sequencer_D1457 =  pf_vf_mux_system_env_TB4_D2.master[107].sequencer;   
    sequencer.master_sequencer_D1458 =  pf_vf_mux_system_env_TB4_D2.master[108].sequencer;   
    sequencer.master_sequencer_D1459 =  pf_vf_mux_system_env_TB4_D2.master[109].sequencer;   
    sequencer.master_sequencer_D1460 =  pf_vf_mux_system_env_TB4_D2.master[110].sequencer;   
    sequencer.master_sequencer_D1461 =  pf_vf_mux_system_env_TB4_D2.master[111].sequencer;   
    sequencer.master_sequencer_D1462 =  pf_vf_mux_system_env_TB4_D2.master[112].sequencer;   
    sequencer.master_sequencer_D1463 =  pf_vf_mux_system_env_TB4_D2.master[113].sequencer;   
    sequencer.master_sequencer_D1464 =  pf_vf_mux_system_env_TB4_D2.master[114].sequencer;   
    sequencer.master_sequencer_D1465 =  pf_vf_mux_system_env_TB4_D2.master[115].sequencer;   
    sequencer.master_sequencer_D1466 =  pf_vf_mux_system_env_TB4_D2.master[116].sequencer;   
    sequencer.master_sequencer_D1467 =  pf_vf_mux_system_env_TB4_D2.master[117].sequencer;   
    sequencer.master_sequencer_D1468 =  pf_vf_mux_system_env_TB4_D2.master[118].sequencer;   
    sequencer.master_sequencer_D1469 =  pf_vf_mux_system_env_TB4_D2.master[119].sequencer;   
    sequencer.master_sequencer_D1470 =  pf_vf_mux_system_env_TB4_D2.master[120].sequencer;   
    sequencer.master_sequencer_D1471 =  pf_vf_mux_system_env_TB4_D2.master[121].sequencer;   
    sequencer.master_sequencer_D1472 =  pf_vf_mux_system_env_TB4_D2.master[122].sequencer;   
    sequencer.master_sequencer_D1473 =  pf_vf_mux_system_env_TB4_D2.master[123].sequencer;   
    sequencer.master_sequencer_D1474 =  pf_vf_mux_system_env_TB4_D2.master[124].sequencer;   
    sequencer.master_sequencer_D1475 =  pf_vf_mux_system_env_TB4_D2.master[125].sequencer;   
    sequencer.master_sequencer_D1476 =  pf_vf_mux_system_env_TB4_D2.master[126].sequencer;   
    sequencer.master_sequencer_D1477 =  pf_vf_mux_system_env_TB4_D2.master[127].sequencer;   
    sequencer.master_sequencer_D1478 =  pf_vf_mux_system_env_TB4_D2.master[128].sequencer;   
    sequencer.master_sequencer_D1479 =  pf_vf_mux_system_env_TB4_D2.master[129].sequencer;   
    sequencer.master_sequencer_D1480 =  pf_vf_mux_system_env_TB4_D2.master[130].sequencer;   
    sequencer.master_sequencer_D1481 =  pf_vf_mux_system_env_TB4_D2.master[131].sequencer;   
    sequencer.master_sequencer_D1482 =  pf_vf_mux_system_env_TB4_D2.master[132].sequencer;   
    sequencer.master_sequencer_D1483 =  pf_vf_mux_system_env_TB4_D2.master[133].sequencer;   
    sequencer.master_sequencer_D1484 =  pf_vf_mux_system_env_TB4_D2.master[134].sequencer;   
    sequencer.master_sequencer_D1485 =  pf_vf_mux_system_env_TB4_D2.master[135].sequencer;   
    sequencer.master_sequencer_D1486 =  pf_vf_mux_system_env_TB4_D2.master[136].sequencer;   
    sequencer.master_sequencer_D1487 =  pf_vf_mux_system_env_TB4_D2.master[137].sequencer;   
    sequencer.master_sequencer_D1488 =  pf_vf_mux_system_env_TB4_D2.master[138].sequencer;   
    sequencer.master_sequencer_D1489 =  pf_vf_mux_system_env_TB4_D2.master[139].sequencer;   
    sequencer.master_sequencer_D1490 =  pf_vf_mux_system_env_TB4_D2.master[140].sequencer;   
    sequencer.master_sequencer_D1491 =  pf_vf_mux_system_env_TB4_D2.master[141].sequencer;   
    sequencer.master_sequencer_D1492 =  pf_vf_mux_system_env_TB4_D2.master[142].sequencer;   
    sequencer.master_sequencer_D1493 =  pf_vf_mux_system_env_TB4_D2.master[143].sequencer;   
    sequencer.master_sequencer_D1494 =  pf_vf_mux_system_env_TB4_D2.master[144].sequencer;   
    sequencer.master_sequencer_D1495 =  pf_vf_mux_system_env_TB4_D2.master[145].sequencer;   
    sequencer.master_sequencer_D1496 =  pf_vf_mux_system_env_TB4_D2.master[146].sequencer;   
    sequencer.master_sequencer_D1497 =  pf_vf_mux_system_env_TB4_D2.master[147].sequencer;   
    sequencer.master_sequencer_D1498 =  pf_vf_mux_system_env_TB4_D2.master[148].sequencer;   
    sequencer.master_sequencer_D1499 =  pf_vf_mux_system_env_TB4_D2.master[149].sequencer;   
    sequencer.master_sequencer_D1500 =  pf_vf_mux_system_env_TB4_D2.master[150].sequencer;   
    sequencer.master_sequencer_D1501 =  pf_vf_mux_system_env_TB4_D2.master[151].sequencer;   
    sequencer.master_sequencer_D1502 =  pf_vf_mux_system_env_TB4_D2.master[152].sequencer;   
    sequencer.master_sequencer_D1503 =  pf_vf_mux_system_env_TB4_D2.master[153].sequencer;   
    sequencer.master_sequencer_D1504 =  pf_vf_mux_system_env_TB4_D2.master[154].sequencer;   
    sequencer.master_sequencer_D1505 =  pf_vf_mux_system_env_TB4_D2.master[155].sequencer;   
    sequencer.master_sequencer_D1506 =  pf_vf_mux_system_env_TB4_D2.master[156].sequencer;   
    sequencer.master_sequencer_D1507 =  pf_vf_mux_system_env_TB4_D2.master[157].sequencer;   
    sequencer.master_sequencer_D1508 =  pf_vf_mux_system_env_TB4_D2.master[158].sequencer;   
    sequencer.master_sequencer_D1509 =  pf_vf_mux_system_env_TB4_D2.master[159].sequencer;   
    sequencer.master_sequencer_D1510 =  pf_vf_mux_system_env_TB4_D2.master[160].sequencer;   
    sequencer.master_sequencer_D1511 =  pf_vf_mux_system_env_TB4_D2.master[161].sequencer;   
    sequencer.master_sequencer_D1512 =  pf_vf_mux_system_env_TB4_D2.master[162].sequencer;   
    sequencer.master_sequencer_D1513 =  pf_vf_mux_system_env_TB4_D2.master[163].sequencer;   
    sequencer.master_sequencer_D1514 =  pf_vf_mux_system_env_TB4_D2.master[164].sequencer;   
    sequencer.master_sequencer_D1515 =  pf_vf_mux_system_env_TB4_D2.master[165].sequencer;   
    sequencer.master_sequencer_D1516 =  pf_vf_mux_system_env_TB4_D2.master[166].sequencer;   
    sequencer.master_sequencer_D1517 =  pf_vf_mux_system_env_TB4_D2.master[167].sequencer;   
    sequencer.master_sequencer_D1518 =  pf_vf_mux_system_env_TB4_D2.master[168].sequencer;   
    sequencer.master_sequencer_D1519 =  pf_vf_mux_system_env_TB4_D2.master[169].sequencer;   
    sequencer.master_sequencer_D1520 =  pf_vf_mux_system_env_TB4_D2.master[170].sequencer;   
    sequencer.master_sequencer_D1521 =  pf_vf_mux_system_env_TB4_D2.master[171].sequencer;   
    sequencer.master_sequencer_D1522 =  pf_vf_mux_system_env_TB4_D2.master[172].sequencer;   
    sequencer.master_sequencer_D1523 =  pf_vf_mux_system_env_TB4_D2.master[173].sequencer;   
    sequencer.master_sequencer_D1524 =  pf_vf_mux_system_env_TB4_D2.master[174].sequencer;   
    sequencer.master_sequencer_D1525 =  pf_vf_mux_system_env_TB4_D2.master[175].sequencer;   
    sequencer.master_sequencer_D1526 =  pf_vf_mux_system_env_TB4_D2.master[176].sequencer;   
    sequencer.master_sequencer_D1527 =  pf_vf_mux_system_env_TB4_D2.master[177].sequencer;   
    sequencer.master_sequencer_D1528 =  pf_vf_mux_system_env_TB4_D2.master[178].sequencer;   
    sequencer.master_sequencer_D1529 =  pf_vf_mux_system_env_TB4_D2.master[179].sequencer;   
    sequencer.master_sequencer_D1530 =  pf_vf_mux_system_env_TB4_D2.master[180].sequencer;   
    sequencer.master_sequencer_D1531 =  pf_vf_mux_system_env_TB4_D2.master[181].sequencer;   
    sequencer.master_sequencer_D1532 =  pf_vf_mux_system_env_TB4_D2.master[182].sequencer;   
    sequencer.master_sequencer_D1533 =  pf_vf_mux_system_env_TB4_D2.master[183].sequencer;   
    sequencer.master_sequencer_D1534 =  pf_vf_mux_system_env_TB4_D2.master[184].sequencer;   
    sequencer.master_sequencer_D1535 =  pf_vf_mux_system_env_TB4_D2.master[185].sequencer;   
    sequencer.master_sequencer_D1536 =  pf_vf_mux_system_env_TB4_D2.master[186].sequencer;   
    sequencer.master_sequencer_D1537 =  pf_vf_mux_system_env_TB4_D2.master[187].sequencer;   
    sequencer.master_sequencer_D1538 =  pf_vf_mux_system_env_TB4_D2.master[188].sequencer;   
    sequencer.master_sequencer_D1539 =  pf_vf_mux_system_env_TB4_D2.master[189].sequencer;   
    sequencer.master_sequencer_D1540 =  pf_vf_mux_system_env_TB4_D2.master[190].sequencer;   
    sequencer.master_sequencer_D1541 =  pf_vf_mux_system_env_TB4_D2.master[191].sequencer;   
    sequencer.master_sequencer_D1542 =  pf_vf_mux_system_env_TB4_D2.master[192].sequencer;   
    sequencer.master_sequencer_D1543 =  pf_vf_mux_system_env_TB4_D2.master[193].sequencer;   
    sequencer.master_sequencer_D1544 =  pf_vf_mux_system_env_TB4_D2.master[194].sequencer;   
    sequencer.master_sequencer_D1545 =  pf_vf_mux_system_env_TB4_D2.master[195].sequencer;   
    sequencer.master_sequencer_D1546 =  pf_vf_mux_system_env_TB4_D2.master[196].sequencer;   
    sequencer.master_sequencer_D1547 =  pf_vf_mux_system_env_TB4_D2.master[197].sequencer;   
    sequencer.master_sequencer_D1548 =  pf_vf_mux_system_env_TB4_D2.master[198].sequencer;   
    sequencer.master_sequencer_D1549 =  pf_vf_mux_system_env_TB4_D2.master[199].sequencer;   
    sequencer.master_sequencer_D1550 =  pf_vf_mux_system_env_TB4_D2.master[200].sequencer;   
    sequencer.master_sequencer_D1551 =  pf_vf_mux_system_env_TB4_D2.master[201].sequencer;   
    sequencer.master_sequencer_D1552 =  pf_vf_mux_system_env_TB4_D2.master[202].sequencer;   
    sequencer.master_sequencer_D1553 =  pf_vf_mux_system_env_TB4_D2.master[203].sequencer;   
    sequencer.master_sequencer_D1554 =  pf_vf_mux_system_env_TB4_D2.master[204].sequencer;   
    sequencer.master_sequencer_D1555 =  pf_vf_mux_system_env_TB4_D2.master[205].sequencer;   
    sequencer.master_sequencer_D1556 =  pf_vf_mux_system_env_TB4_D2.master[206].sequencer;   
    sequencer.master_sequencer_D1557 =  pf_vf_mux_system_env_TB4_D2.master[207].sequencer;   
    sequencer.master_sequencer_D1558 =  pf_vf_mux_system_env_TB4_D2.master[208].sequencer;   
    sequencer.master_sequencer_D1559 =  pf_vf_mux_system_env_TB4_D2.master[209].sequencer;   
    sequencer.master_sequencer_D1560 =  pf_vf_mux_system_env_TB4_D2.master[210].sequencer;   
    sequencer.master_sequencer_D1561 =  pf_vf_mux_system_env_TB4_D2.master[211].sequencer;   
    sequencer.master_sequencer_D1562 =  pf_vf_mux_system_env_TB4_D2.master[212].sequencer;   
    sequencer.master_sequencer_D1563 =  pf_vf_mux_system_env_TB4_D2.master[213].sequencer;   
    sequencer.master_sequencer_D1564 =  pf_vf_mux_system_env_TB4_D2.master[214].sequencer;   
    sequencer.master_sequencer_D1565 =  pf_vf_mux_system_env_TB4_D2.master[215].sequencer;   
    sequencer.master_sequencer_D1566 =  pf_vf_mux_system_env_TB4_D2.master[216].sequencer;   
    sequencer.master_sequencer_D1567 =  pf_vf_mux_system_env_TB4_D2.master[217].sequencer;   
    sequencer.master_sequencer_D1568 =  pf_vf_mux_system_env_TB4_D2.master[218].sequencer;   
    sequencer.master_sequencer_D1569 =  pf_vf_mux_system_env_TB4_D2.master[219].sequencer;   
    sequencer.master_sequencer_D1570 =  pf_vf_mux_system_env_TB4_D2.master[220].sequencer;   
    sequencer.master_sequencer_D1571 =  pf_vf_mux_system_env_TB4_D2.master[221].sequencer;   
    sequencer.master_sequencer_D1572 =  pf_vf_mux_system_env_TB4_D2.master[222].sequencer;   
    sequencer.master_sequencer_D1573 =  pf_vf_mux_system_env_TB4_D2.master[223].sequencer;   
    sequencer.master_sequencer_D1574 =  pf_vf_mux_system_env_TB4_D2.master[224].sequencer;   
    sequencer.master_sequencer_D1575 =  pf_vf_mux_system_env_TB4_D2.master[225].sequencer;   
    sequencer.master_sequencer_D1576 =  pf_vf_mux_system_env_TB4_D2.master[226].sequencer;   
    sequencer.master_sequencer_D1577 =  pf_vf_mux_system_env_TB4_D2.master[227].sequencer;   
    sequencer.master_sequencer_D1578 =  pf_vf_mux_system_env_TB4_D2.master[228].sequencer;   
    sequencer.master_sequencer_D1579 =  pf_vf_mux_system_env_TB4_D2.master[229].sequencer;   
    sequencer.master_sequencer_D1580 =  pf_vf_mux_system_env_TB4_D2.master[230].sequencer;   
    sequencer.master_sequencer_D1581 =  pf_vf_mux_system_env_TB4_D2.master[231].sequencer;   
    sequencer.master_sequencer_D1582 =  pf_vf_mux_system_env_TB4_D2.master[232].sequencer;   
    sequencer.master_sequencer_D1583 =  pf_vf_mux_system_env_TB4_D2.master[233].sequencer;   
    sequencer.master_sequencer_D1584 =  pf_vf_mux_system_env_TB4_D2.master[234].sequencer;   
    sequencer.master_sequencer_D1585 =  pf_vf_mux_system_env_TB4_D2.master[235].sequencer;   
    sequencer.master_sequencer_D1586 =  pf_vf_mux_system_env_TB4_D2.master[236].sequencer;   
    sequencer.master_sequencer_D1587 =  pf_vf_mux_system_env_TB4_D2.master[237].sequencer;   
    sequencer.master_sequencer_D1588 =  pf_vf_mux_system_env_TB4_D2.master[238].sequencer;   
    sequencer.master_sequencer_D1589 =  pf_vf_mux_system_env_TB4_D2.master[239].sequencer;   
    sequencer.master_sequencer_D1590 =  pf_vf_mux_system_env_TB4_D2.master[240].sequencer;   
    sequencer.master_sequencer_D1591 =  pf_vf_mux_system_env_TB4_D2.master[241].sequencer;   
    sequencer.master_sequencer_D1592 =  pf_vf_mux_system_env_TB4_D2.master[242].sequencer;   
    sequencer.master_sequencer_D1593 =  pf_vf_mux_system_env_TB4_D2.master[243].sequencer;   
    sequencer.master_sequencer_D1594 =  pf_vf_mux_system_env_TB4_D2.master[244].sequencer;   
    sequencer.master_sequencer_D1595 =  pf_vf_mux_system_env_TB4_D2.master[245].sequencer;   
    sequencer.master_sequencer_D1596 =  pf_vf_mux_system_env_TB4_D2.master[246].sequencer;   
    sequencer.master_sequencer_D1597 =  pf_vf_mux_system_env_TB4_D2.master[247].sequencer;   
    sequencer.master_sequencer_D1598 =  pf_vf_mux_system_env_TB4_D2.master[248].sequencer;   
    sequencer.master_sequencer_D1599 =  pf_vf_mux_system_env_TB4_D2.master[249].sequencer;   
    sequencer.master_sequencer_D1600 =  pf_vf_mux_system_env_TB4_D2.master[250].sequencer;   
    sequencer.master_sequencer_D1601 =  pf_vf_mux_system_env_TB4_D2.master[251].sequencer;   
    sequencer.master_sequencer_D1602 =  pf_vf_mux_system_env_TB4_D2.master[252].sequencer;   
    sequencer.master_sequencer_D1603 =  pf_vf_mux_system_env_TB4_D2.master[253].sequencer;   
    sequencer.master_sequencer_D1604 =  pf_vf_mux_system_env_TB4_D2.master[254].sequencer;   
    sequencer.master_sequencer_D1605 =  pf_vf_mux_system_env_TB4_D2.master[255].sequencer;   
    sequencer.master_sequencer_D1606 =  pf_vf_mux_system_env_TB4_D2.master[256].sequencer;   
    sequencer.master_sequencer_D1607 =  pf_vf_mux_system_env_TB4_D2.master[257].sequencer;   
    sequencer.master_sequencer_D1608 =  pf_vf_mux_system_env_TB4_D2.master[258].sequencer;   
    sequencer.master_sequencer_D1609 =  pf_vf_mux_system_env_TB4_D2.master[259].sequencer;   
    sequencer.master_sequencer_D1610 =  pf_vf_mux_system_env_TB4_D2.master[260].sequencer;   
    sequencer.master_sequencer_D1611 =  pf_vf_mux_system_env_TB4_D2.master[261].sequencer;   
    sequencer.master_sequencer_D1612 =  pf_vf_mux_system_env_TB4_D2.master[262].sequencer;   
    sequencer.master_sequencer_D1613 =  pf_vf_mux_system_env_TB4_D2.master[263].sequencer;   
    sequencer.master_sequencer_D1614 =  pf_vf_mux_system_env_TB4_D2.master[264].sequencer;   
    sequencer.master_sequencer_D1615 =  pf_vf_mux_system_env_TB4_D2.master[265].sequencer;   
    sequencer.master_sequencer_D1616 =  pf_vf_mux_system_env_TB4_D2.master[266].sequencer;   
    sequencer.master_sequencer_D1617 =  pf_vf_mux_system_env_TB4_D2.master[267].sequencer;   
    sequencer.master_sequencer_D1618 =  pf_vf_mux_system_env_TB4_D2.master[268].sequencer;   
    sequencer.master_sequencer_D1619 =  pf_vf_mux_system_env_TB4_D2.master[269].sequencer;   
    sequencer.master_sequencer_D1620 =  pf_vf_mux_system_env_TB4_D2.master[270].sequencer;   
    sequencer.master_sequencer_D1621 =  pf_vf_mux_system_env_TB4_D2.master[271].sequencer;   
    sequencer.master_sequencer_D1622 =  pf_vf_mux_system_env_TB4_D2.master[272].sequencer;   
    sequencer.master_sequencer_D1623 =  pf_vf_mux_system_env_TB4_D2.master[273].sequencer;   
    sequencer.master_sequencer_D1624 =  pf_vf_mux_system_env_TB4_D2.master[274].sequencer;   
    sequencer.master_sequencer_D1625 =  pf_vf_mux_system_env_TB4_D2.master[275].sequencer;   
    sequencer.master_sequencer_D1626 =  pf_vf_mux_system_env_TB4_D2.master[276].sequencer;   
    sequencer.master_sequencer_D1627 =  pf_vf_mux_system_env_TB4_D2.master[277].sequencer;   
    sequencer.master_sequencer_D1628 =  pf_vf_mux_system_env_TB4_D2.master[278].sequencer;   
    sequencer.master_sequencer_D1629 =  pf_vf_mux_system_env_TB4_D2.master[279].sequencer;   
    sequencer.master_sequencer_D1630 =  pf_vf_mux_system_env_TB4_D2.master[280].sequencer;   
    sequencer.master_sequencer_D1631 =  pf_vf_mux_system_env_TB4_D2.master[281].sequencer;   
    sequencer.master_sequencer_D1632 =  pf_vf_mux_system_env_TB4_D2.master[282].sequencer;   
    sequencer.master_sequencer_D1633 =  pf_vf_mux_system_env_TB4_D2.master[283].sequencer;   
    sequencer.master_sequencer_D1634 =  pf_vf_mux_system_env_TB4_D2.master[284].sequencer;   
    sequencer.master_sequencer_D1635 =  pf_vf_mux_system_env_TB4_D2.master[285].sequencer;   
    sequencer.master_sequencer_D1636 =  pf_vf_mux_system_env_TB4_D2.master[286].sequencer;   
    sequencer.master_sequencer_D1637 =  pf_vf_mux_system_env_TB4_D2.master[287].sequencer;   
    sequencer.master_sequencer_D1638 =  pf_vf_mux_system_env_TB4_D2.master[288].sequencer;   
    sequencer.master_sequencer_D1639 =  pf_vf_mux_system_env_TB4_D2.master[289].sequencer;   
    sequencer.master_sequencer_D1640 =  pf_vf_mux_system_env_TB4_D2.master[290].sequencer;   
    sequencer.master_sequencer_D1641 =  pf_vf_mux_system_env_TB4_D2.master[291].sequencer;   
    sequencer.master_sequencer_D1642 =  pf_vf_mux_system_env_TB4_D2.master[292].sequencer;   
    sequencer.master_sequencer_D1643 =  pf_vf_mux_system_env_TB4_D2.master[293].sequencer;   
    sequencer.master_sequencer_D1644 =  pf_vf_mux_system_env_TB4_D2.master[294].sequencer;   
    sequencer.master_sequencer_D1645 =  pf_vf_mux_system_env_TB4_D2.master[295].sequencer;   
    sequencer.master_sequencer_D1646 =  pf_vf_mux_system_env_TB4_D2.master[296].sequencer;   
    sequencer.master_sequencer_D1647 =  pf_vf_mux_system_env_TB4_D2.master[297].sequencer;   
    sequencer.master_sequencer_D1648 =  pf_vf_mux_system_env_TB4_D2.master[298].sequencer;   
    sequencer.master_sequencer_D1649 =  pf_vf_mux_system_env_TB4_D2.master[299].sequencer;   
    sequencer.master_sequencer_D1650 =  pf_vf_mux_system_env_TB4_D2.master[300].sequencer;   
    sequencer.master_sequencer_D1651 =  pf_vf_mux_system_env_TB4_D2.master[301].sequencer;   
    sequencer.master_sequencer_D1652 =  pf_vf_mux_system_env_TB4_D2.master[302].sequencer;   
    sequencer.master_sequencer_D1653 =  pf_vf_mux_system_env_TB4_D2.master[303].sequencer;   
    sequencer.master_sequencer_D1654 =  pf_vf_mux_system_env_TB4_D2.master[304].sequencer;   
    sequencer.master_sequencer_D1655 =  pf_vf_mux_system_env_TB4_D2.master[305].sequencer;   
    sequencer.master_sequencer_D1656 =  pf_vf_mux_system_env_TB4_D2.master[306].sequencer;   
    sequencer.master_sequencer_D1657 =  pf_vf_mux_system_env_TB4_D2.master[307].sequencer;   
    sequencer.master_sequencer_D1658 =  pf_vf_mux_system_env_TB4_D2.master[308].sequencer;   
    sequencer.master_sequencer_D1659 =  pf_vf_mux_system_env_TB4_D2.master[309].sequencer;   
    sequencer.master_sequencer_D1660 =  pf_vf_mux_system_env_TB4_D2.master[310].sequencer;   
    sequencer.master_sequencer_D1661 =  pf_vf_mux_system_env_TB4_D2.master[311].sequencer;   
    sequencer.master_sequencer_D1662 =  pf_vf_mux_system_env_TB4_D2.master[312].sequencer;   
    sequencer.master_sequencer_D1663 =  pf_vf_mux_system_env_TB4_D2.master[313].sequencer;   
    sequencer.master_sequencer_D1664 =  pf_vf_mux_system_env_TB4_D2.master[314].sequencer;   
    sequencer.master_sequencer_D1665 =  pf_vf_mux_system_env_TB4_D2.master[315].sequencer;   
    sequencer.master_sequencer_D1666 =  pf_vf_mux_system_env_TB4_D2.master[316].sequencer;   
    sequencer.master_sequencer_D1667 =  pf_vf_mux_system_env_TB4_D2.master[317].sequencer;   
    sequencer.master_sequencer_D1668 =  pf_vf_mux_system_env_TB4_D2.master[318].sequencer;   
    sequencer.master_sequencer_D1669 =  pf_vf_mux_system_env_TB4_D2.master[319].sequencer;   
    sequencer.master_sequencer_D1670 =  pf_vf_mux_system_env_TB4_D2.master[320].sequencer;   
    sequencer.master_sequencer_D1671 =  pf_vf_mux_system_env_TB4_D2.master[321].sequencer;   
    sequencer.master_sequencer_D1672 =  pf_vf_mux_system_env_TB4_D2.master[322].sequencer;   
    sequencer.master_sequencer_D1673 =  pf_vf_mux_system_env_TB4_D2.master[323].sequencer;   
    sequencer.master_sequencer_D1674 =  pf_vf_mux_system_env_TB4_D2.master[324].sequencer;   
    sequencer.master_sequencer_D1675 =  pf_vf_mux_system_env_TB4_D2.master[325].sequencer;   
    sequencer.master_sequencer_D1676 =  pf_vf_mux_system_env_TB4_D2.master[326].sequencer;   
    sequencer.master_sequencer_D1677 =  pf_vf_mux_system_env_TB4_D2.master[327].sequencer;   
    sequencer.master_sequencer_D1678 =  pf_vf_mux_system_env_TB4_D2.master[328].sequencer;   
    sequencer.master_sequencer_D1679 =  pf_vf_mux_system_env_TB4_D2.master[329].sequencer;   
    sequencer.master_sequencer_D1680 =  pf_vf_mux_system_env_TB4_D2.master[330].sequencer;   
    sequencer.master_sequencer_D1681 =  pf_vf_mux_system_env_TB4_D2.master[331].sequencer;   
    sequencer.master_sequencer_D1682 =  pf_vf_mux_system_env_TB4_D2.master[332].sequencer;   
    sequencer.master_sequencer_D1683 =  pf_vf_mux_system_env_TB4_D2.master[333].sequencer;   
    sequencer.master_sequencer_D1684 =  pf_vf_mux_system_env_TB4_D2.master[334].sequencer;   
    sequencer.master_sequencer_D1685 =  pf_vf_mux_system_env_TB4_D2.master[335].sequencer;   
    sequencer.master_sequencer_D1686 =  pf_vf_mux_system_env_TB4_D2.master[336].sequencer;   
    sequencer.master_sequencer_D1687 =  pf_vf_mux_system_env_TB4_D2.master[337].sequencer;   
    sequencer.master_sequencer_D1688 =  pf_vf_mux_system_env_TB4_D2.master[338].sequencer;   
    sequencer.master_sequencer_D1689 =  pf_vf_mux_system_env_TB4_D2.master[339].sequencer;   
    sequencer.master_sequencer_D1690 =  pf_vf_mux_system_env_TB4_D2.master[340].sequencer;   
    sequencer.master_sequencer_D1691 =  pf_vf_mux_system_env_TB4_D2.master[341].sequencer;   
    sequencer.master_sequencer_D1692 =  pf_vf_mux_system_env_TB4_D2.master[342].sequencer;   
    sequencer.master_sequencer_D1693 =  pf_vf_mux_system_env_TB4_D2.master[343].sequencer;   
    sequencer.master_sequencer_D1694 =  pf_vf_mux_system_env_TB4_D2.master[344].sequencer;   
    sequencer.master_sequencer_D1695 =  pf_vf_mux_system_env_TB4_D2.master[345].sequencer;   
    sequencer.master_sequencer_D1696 =  pf_vf_mux_system_env_TB4_D2.master[346].sequencer;   
    sequencer.master_sequencer_D1697 =  pf_vf_mux_system_env_TB4_D2.master[347].sequencer;   
    sequencer.master_sequencer_D1698 =  pf_vf_mux_system_env_TB4_D2.master[348].sequencer;   
    sequencer.master_sequencer_D1699 =  pf_vf_mux_system_env_TB4_D2.master[349].sequencer;   
    sequencer.master_sequencer_D1700 =  pf_vf_mux_system_env_TB4_D2.master[350].sequencer;   
    sequencer.master_sequencer_D1701 =  pf_vf_mux_system_env_TB4_D2.master[351].sequencer;   
    sequencer.master_sequencer_D1702 =  pf_vf_mux_system_env_TB4_D2.master[352].sequencer;   
    sequencer.master_sequencer_D1703 =  pf_vf_mux_system_env_TB4_D2.master[353].sequencer;   
    sequencer.master_sequencer_D1704 =  pf_vf_mux_system_env_TB4_D2.master[354].sequencer;   
    sequencer.master_sequencer_D1705 =  pf_vf_mux_system_env_TB4_D2.master[355].sequencer;   
    sequencer.master_sequencer_D1706 =  pf_vf_mux_system_env_TB4_D2.master[356].sequencer;   
    sequencer.master_sequencer_D1707 =  pf_vf_mux_system_env_TB4_D2.master[357].sequencer;   
    sequencer.master_sequencer_D1708 =  pf_vf_mux_system_env_TB4_D2.master[358].sequencer;   
    sequencer.master_sequencer_D1709 =  pf_vf_mux_system_env_TB4_D2.master[359].sequencer;   
    sequencer.master_sequencer_D1710 =  pf_vf_mux_system_env_TB4_D2.master[360].sequencer;   
    sequencer.master_sequencer_D1711 =  pf_vf_mux_system_env_TB4_D2.master[361].sequencer;   
    sequencer.master_sequencer_D1712 =  pf_vf_mux_system_env_TB4_D2.master[362].sequencer;   
    sequencer.master_sequencer_D1713 =  pf_vf_mux_system_env_TB4_D2.master[363].sequencer;   
    sequencer.master_sequencer_D1714 =  pf_vf_mux_system_env_TB4_D2.master[364].sequencer;   
    sequencer.master_sequencer_D1715 =  pf_vf_mux_system_env_TB4_D2.master[365].sequencer;   
    sequencer.master_sequencer_D1716 =  pf_vf_mux_system_env_TB4_D2.master[366].sequencer;   
    sequencer.master_sequencer_D1717 =  pf_vf_mux_system_env_TB4_D2.master[367].sequencer;   
    sequencer.master_sequencer_D1718 =  pf_vf_mux_system_env_TB4_D2.master[368].sequencer;   
    sequencer.master_sequencer_D1719 =  pf_vf_mux_system_env_TB4_D2.master[369].sequencer;   
    sequencer.master_sequencer_D1720 =  pf_vf_mux_system_env_TB4_D2.master[370].sequencer;   
    sequencer.master_sequencer_D1721 =  pf_vf_mux_system_env_TB4_D2.master[371].sequencer;   
    sequencer.master_sequencer_D1722 =  pf_vf_mux_system_env_TB4_D2.master[372].sequencer;   
    sequencer.master_sequencer_D1723 =  pf_vf_mux_system_env_TB4_D2.master[373].sequencer;   
    sequencer.master_sequencer_D1724 =  pf_vf_mux_system_env_TB4_D2.master[374].sequencer;   
    sequencer.master_sequencer_D1725 =  pf_vf_mux_system_env_TB4_D2.master[375].sequencer;   
    sequencer.master_sequencer_D1726 =  pf_vf_mux_system_env_TB4_D2.master[376].sequencer;   
    sequencer.master_sequencer_D1727 =  pf_vf_mux_system_env_TB4_D2.master[377].sequencer;   
    sequencer.master_sequencer_D1728 =  pf_vf_mux_system_env_TB4_D2.master[378].sequencer;   
    sequencer.master_sequencer_D1729 =  pf_vf_mux_system_env_TB4_D2.master[379].sequencer;   
    sequencer.master_sequencer_D1730 =  pf_vf_mux_system_env_TB4_D2.master[380].sequencer;   
    sequencer.master_sequencer_D1731 =  pf_vf_mux_system_env_TB4_D2.master[381].sequencer;   
    sequencer.master_sequencer_D1732 =  pf_vf_mux_system_env_TB4_D2.master[382].sequencer;   
    sequencer.master_sequencer_D1733 =  pf_vf_mux_system_env_TB4_D2.master[383].sequencer;   
    sequencer.master_sequencer_D1734 =  pf_vf_mux_system_env_TB4_D2.master[384].sequencer;   
    sequencer.master_sequencer_D1735 =  pf_vf_mux_system_env_TB4_D2.master[385].sequencer;   
    sequencer.master_sequencer_D1736 =  pf_vf_mux_system_env_TB4_D2.master[386].sequencer;   
    sequencer.master_sequencer_D1737 =  pf_vf_mux_system_env_TB4_D2.master[387].sequencer;   
    sequencer.master_sequencer_D1738 =  pf_vf_mux_system_env_TB4_D2.master[388].sequencer;   
    sequencer.master_sequencer_D1739 =  pf_vf_mux_system_env_TB4_D2.master[389].sequencer;   
    sequencer.master_sequencer_D1740 =  pf_vf_mux_system_env_TB4_D2.master[390].sequencer;   
    sequencer.master_sequencer_D1741 =  pf_vf_mux_system_env_TB4_D2.master[391].sequencer;   
    sequencer.master_sequencer_D1742 =  pf_vf_mux_system_env_TB4_D2.master[392].sequencer;   
    sequencer.master_sequencer_D1743 =  pf_vf_mux_system_env_TB4_D2.master[393].sequencer;   
    sequencer.master_sequencer_D1744 =  pf_vf_mux_system_env_TB4_D2.master[394].sequencer;   
    sequencer.master_sequencer_D1745 =  pf_vf_mux_system_env_TB4_D2.master[395].sequencer;   
    sequencer.master_sequencer_D1746 =  pf_vf_mux_system_env_TB4_D2.master[396].sequencer;   
    sequencer.master_sequencer_D1747 =  pf_vf_mux_system_env_TB4_D2.master[397].sequencer;   
    sequencer.master_sequencer_D1748 =  pf_vf_mux_system_env_TB4_D2.master[398].sequencer;   
    sequencer.master_sequencer_D1749 =  pf_vf_mux_system_env_TB4_D2.master[399].sequencer;   
    sequencer.master_sequencer_D1750 =  pf_vf_mux_system_env_TB4_D2.master[400].sequencer;   
    sequencer.master_sequencer_D1751 =  pf_vf_mux_system_env_TB4_D2.master[401].sequencer;   
    sequencer.master_sequencer_D1752 =  pf_vf_mux_system_env_TB4_D2.master[402].sequencer;   
    sequencer.master_sequencer_D1753 =  pf_vf_mux_system_env_TB4_D2.master[403].sequencer;   
    sequencer.master_sequencer_D1754 =  pf_vf_mux_system_env_TB4_D2.master[404].sequencer;   
    sequencer.master_sequencer_D1755 =  pf_vf_mux_system_env_TB4_D2.master[405].sequencer;   
    sequencer.master_sequencer_D1756 =  pf_vf_mux_system_env_TB4_D2.master[406].sequencer;   
    sequencer.master_sequencer_D1757 =  pf_vf_mux_system_env_TB4_D2.master[407].sequencer;   
    sequencer.master_sequencer_D1758 =  pf_vf_mux_system_env_TB4_D2.master[408].sequencer;   
    sequencer.master_sequencer_D1759 =  pf_vf_mux_system_env_TB4_D2.master[409].sequencer;   
    sequencer.master_sequencer_D1760 =  pf_vf_mux_system_env_TB4_D2.master[410].sequencer;   
    sequencer.master_sequencer_D1761 =  pf_vf_mux_system_env_TB4_D2.master[411].sequencer;   
    sequencer.master_sequencer_D1762 =  pf_vf_mux_system_env_TB4_D2.master[412].sequencer;   
    sequencer.master_sequencer_D1763 =  pf_vf_mux_system_env_TB4_D2.master[413].sequencer;   
    sequencer.master_sequencer_D1764 =  pf_vf_mux_system_env_TB4_D2.master[414].sequencer;   
    sequencer.master_sequencer_D1765 =  pf_vf_mux_system_env_TB4_D2.master[415].sequencer;   
    sequencer.master_sequencer_D1766 =  pf_vf_mux_system_env_TB4_D2.master[416].sequencer;   
    sequencer.master_sequencer_D1767 =  pf_vf_mux_system_env_TB4_D2.master[417].sequencer;   
    sequencer.master_sequencer_D1768 =  pf_vf_mux_system_env_TB4_D2.master[418].sequencer;   
    sequencer.master_sequencer_D1769 =  pf_vf_mux_system_env_TB4_D2.master[419].sequencer;   
    sequencer.master_sequencer_D1770 =  pf_vf_mux_system_env_TB4_D2.master[420].sequencer;   
    sequencer.master_sequencer_D1771 =  pf_vf_mux_system_env_TB4_D2.master[421].sequencer;   
    sequencer.master_sequencer_D1772 =  pf_vf_mux_system_env_TB4_D2.master[422].sequencer;   
    sequencer.master_sequencer_D1773 =  pf_vf_mux_system_env_TB4_D2.master[423].sequencer;   
    sequencer.master_sequencer_D1774 =  pf_vf_mux_system_env_TB4_D2.master[424].sequencer;   
    sequencer.master_sequencer_D1775 =  pf_vf_mux_system_env_TB4_D2.master[425].sequencer;   
    sequencer.master_sequencer_D1776 =  pf_vf_mux_system_env_TB4_D2.master[426].sequencer;   
    sequencer.master_sequencer_D1777 =  pf_vf_mux_system_env_TB4_D2.master[427].sequencer;   
    sequencer.master_sequencer_D1778 =  pf_vf_mux_system_env_TB4_D2.master[428].sequencer;   
    sequencer.master_sequencer_D1779 =  pf_vf_mux_system_env_TB4_D2.master[429].sequencer;   
    sequencer.master_sequencer_D1780 =  pf_vf_mux_system_env_TB4_D2.master[430].sequencer;   
    sequencer.master_sequencer_D1781 =  pf_vf_mux_system_env_TB4_D2.master[431].sequencer;   
    sequencer.master_sequencer_D1782 =  pf_vf_mux_system_env_TB4_D2.master[432].sequencer;   
    sequencer.master_sequencer_D1783 =  pf_vf_mux_system_env_TB4_D2.master[433].sequencer;   
    sequencer.master_sequencer_D1784 =  pf_vf_mux_system_env_TB4_D2.master[434].sequencer;   
    sequencer.master_sequencer_D1785 =  pf_vf_mux_system_env_TB4_D2.master[435].sequencer;   
    sequencer.master_sequencer_D1786 =  pf_vf_mux_system_env_TB4_D2.master[436].sequencer;   
    sequencer.master_sequencer_D1787 =  pf_vf_mux_system_env_TB4_D2.master[437].sequencer;   
    sequencer.master_sequencer_D1788 =  pf_vf_mux_system_env_TB4_D2.master[438].sequencer;   
    sequencer.master_sequencer_D1789 =  pf_vf_mux_system_env_TB4_D2.master[439].sequencer;   
    sequencer.master_sequencer_D1790 =  pf_vf_mux_system_env_TB4_D2.master[440].sequencer;   
    sequencer.master_sequencer_D1791 =  pf_vf_mux_system_env_TB4_D2.master[441].sequencer;   
    sequencer.master_sequencer_D1792 =  pf_vf_mux_system_env_TB4_D2.master[442].sequencer;   
    sequencer.master_sequencer_D1793 =  pf_vf_mux_system_env_TB4_D2.master[443].sequencer;   
    sequencer.master_sequencer_D1794 =  pf_vf_mux_system_env_TB4_D2.master[444].sequencer;   
    sequencer.master_sequencer_D1795 =  pf_vf_mux_system_env_TB4_D2.master[445].sequencer;   
    sequencer.master_sequencer_D1796 =  pf_vf_mux_system_env_TB4_D2.master[446].sequencer;   
    sequencer.master_sequencer_D1797 =  pf_vf_mux_system_env_TB4_D2.master[447].sequencer;   
    sequencer.master_sequencer_D1798 =  pf_vf_mux_system_env_TB4_D2.master[448].sequencer;   
    sequencer.master_sequencer_D1799 =  pf_vf_mux_system_env_TB4_D2.master[449].sequencer;   
    sequencer.master_sequencer_D1800 =  pf_vf_mux_system_env_TB4_D3.master[0].sequencer;   
    sequencer.master_sequencer_D1801 =  pf_vf_mux_system_env_TB4_D3.master[1].sequencer;   
    sequencer.master_sequencer_D1802 =  pf_vf_mux_system_env_TB4_D3.master[2].sequencer;   
    sequencer.master_sequencer_D1803 =  pf_vf_mux_system_env_TB4_D3.master[3].sequencer;   
    sequencer.master_sequencer_D1804 =  pf_vf_mux_system_env_TB4_D3.master[4].sequencer;   
    sequencer.master_sequencer_D1805 =  pf_vf_mux_system_env_TB4_D3.master[5].sequencer;   
    sequencer.master_sequencer_D1806 =  pf_vf_mux_system_env_TB4_D3.master[6].sequencer;   
    sequencer.master_sequencer_D1807 =  pf_vf_mux_system_env_TB4_D3.master[7].sequencer;   
    sequencer.master_sequencer_D1808 =  pf_vf_mux_system_env_TB4_D3.master[8].sequencer;   
    sequencer.master_sequencer_D1809 =  pf_vf_mux_system_env_TB4_D3.master[9].sequencer;   
    sequencer.master_sequencer_D1810 =  pf_vf_mux_system_env_TB4_D3.master[10].sequencer;   
    sequencer.master_sequencer_D1811 =  pf_vf_mux_system_env_TB4_D3.master[11].sequencer;   
    sequencer.master_sequencer_D1812 =  pf_vf_mux_system_env_TB4_D3.master[12].sequencer;   
    sequencer.master_sequencer_D1813 =  pf_vf_mux_system_env_TB4_D3.master[13].sequencer;   
    sequencer.master_sequencer_D1814 =  pf_vf_mux_system_env_TB4_D3.master[14].sequencer;   
    sequencer.master_sequencer_D1815 =  pf_vf_mux_system_env_TB4_D3.master[15].sequencer;   
    sequencer.master_sequencer_D1816 =  pf_vf_mux_system_env_TB4_D3.master[16].sequencer;   
    sequencer.master_sequencer_D1817 =  pf_vf_mux_system_env_TB4_D3.master[17].sequencer;   
    sequencer.master_sequencer_D1818 =  pf_vf_mux_system_env_TB4_D3.master[18].sequencer;   
    sequencer.master_sequencer_D1819 =  pf_vf_mux_system_env_TB4_D3.master[19].sequencer;   
    sequencer.master_sequencer_D1820 =  pf_vf_mux_system_env_TB4_D3.master[20].sequencer;   
    sequencer.master_sequencer_D1821 =  pf_vf_mux_system_env_TB4_D3.master[21].sequencer;   
    sequencer.master_sequencer_D1822 =  pf_vf_mux_system_env_TB4_D3.master[22].sequencer;   
    sequencer.master_sequencer_D1823 =  pf_vf_mux_system_env_TB4_D3.master[23].sequencer;   
    sequencer.master_sequencer_D1824 =  pf_vf_mux_system_env_TB4_D3.master[24].sequencer;   
    sequencer.master_sequencer_D1825 =  pf_vf_mux_system_env_TB4_D3.master[25].sequencer;   
    sequencer.master_sequencer_D1826 =  pf_vf_mux_system_env_TB4_D3.master[26].sequencer;   
    sequencer.master_sequencer_D1827 =  pf_vf_mux_system_env_TB4_D3.master[27].sequencer;   
    sequencer.master_sequencer_D1828 =  pf_vf_mux_system_env_TB4_D3.master[28].sequencer;   
    sequencer.master_sequencer_D1829 =  pf_vf_mux_system_env_TB4_D3.master[29].sequencer;   
    sequencer.master_sequencer_D1830 =  pf_vf_mux_system_env_TB4_D3.master[30].sequencer;   
    sequencer.master_sequencer_D1831 =  pf_vf_mux_system_env_TB4_D3.master[31].sequencer;   
    sequencer.master_sequencer_D1832 =  pf_vf_mux_system_env_TB4_D3.master[32].sequencer;   
    sequencer.master_sequencer_D1833 =  pf_vf_mux_system_env_TB4_D3.master[33].sequencer;   
    sequencer.master_sequencer_D1834 =  pf_vf_mux_system_env_TB4_D3.master[34].sequencer;   
    sequencer.master_sequencer_D1835 =  pf_vf_mux_system_env_TB4_D3.master[35].sequencer;   
    sequencer.master_sequencer_D1836 =  pf_vf_mux_system_env_TB4_D3.master[36].sequencer;   
    sequencer.master_sequencer_D1837 =  pf_vf_mux_system_env_TB4_D3.master[37].sequencer;   
    sequencer.master_sequencer_D1838 =  pf_vf_mux_system_env_TB4_D3.master[38].sequencer;   
    sequencer.master_sequencer_D1839 =  pf_vf_mux_system_env_TB4_D3.master[39].sequencer;   
    sequencer.master_sequencer_D1840 =  pf_vf_mux_system_env_TB4_D3.master[40].sequencer;   
    sequencer.master_sequencer_D1841 =  pf_vf_mux_system_env_TB4_D3.master[41].sequencer;   
    sequencer.master_sequencer_D1842 =  pf_vf_mux_system_env_TB4_D3.master[42].sequencer;   
    sequencer.master_sequencer_D1843 =  pf_vf_mux_system_env_TB4_D3.master[43].sequencer;   
    sequencer.master_sequencer_D1844 =  pf_vf_mux_system_env_TB4_D3.master[44].sequencer;   
    sequencer.master_sequencer_D1845 =  pf_vf_mux_system_env_TB4_D3.master[45].sequencer;   
    sequencer.master_sequencer_D1846 =  pf_vf_mux_system_env_TB4_D3.master[46].sequencer;   
    sequencer.master_sequencer_D1847 =  pf_vf_mux_system_env_TB4_D3.master[47].sequencer;   
    sequencer.master_sequencer_D1848 =  pf_vf_mux_system_env_TB4_D3.master[48].sequencer;   
    sequencer.master_sequencer_D1849 =  pf_vf_mux_system_env_TB4_D3.master[49].sequencer;   
    sequencer.master_sequencer_D1850 =  pf_vf_mux_system_env_TB4_D3.master[50].sequencer;   
    sequencer.master_sequencer_D1851 =  pf_vf_mux_system_env_TB4_D3.master[51].sequencer;   
    sequencer.master_sequencer_D1852 =  pf_vf_mux_system_env_TB4_D3.master[52].sequencer;   
    sequencer.master_sequencer_D1853 =  pf_vf_mux_system_env_TB4_D3.master[53].sequencer;   
    sequencer.master_sequencer_D1854 =  pf_vf_mux_system_env_TB4_D3.master[54].sequencer;   
    sequencer.master_sequencer_D1855 =  pf_vf_mux_system_env_TB4_D3.master[55].sequencer;   
    sequencer.master_sequencer_D1856 =  pf_vf_mux_system_env_TB4_D3.master[56].sequencer;   
    sequencer.master_sequencer_D1857 =  pf_vf_mux_system_env_TB4_D3.master[57].sequencer;   
    sequencer.master_sequencer_D1858 =  pf_vf_mux_system_env_TB4_D3.master[58].sequencer;   
    sequencer.master_sequencer_D1859 =  pf_vf_mux_system_env_TB4_D3.master[59].sequencer;   
    sequencer.master_sequencer_D1860 =  pf_vf_mux_system_env_TB4_D3.master[60].sequencer;   
    sequencer.master_sequencer_D1861 =  pf_vf_mux_system_env_TB4_D3.master[61].sequencer;   
    sequencer.master_sequencer_D1862 =  pf_vf_mux_system_env_TB4_D3.master[62].sequencer;   
    sequencer.master_sequencer_D1863 =  pf_vf_mux_system_env_TB4_D3.master[63].sequencer;   
    sequencer.master_sequencer_D1864 =  pf_vf_mux_system_env_TB4_D3.master[64].sequencer;   
    sequencer.master_sequencer_D1865 =  pf_vf_mux_system_env_TB4_D3.master[65].sequencer;   
    sequencer.master_sequencer_D1866 =  pf_vf_mux_system_env_TB4_D3.master[66].sequencer;   
    sequencer.master_sequencer_D1867 =  pf_vf_mux_system_env_TB4_D3.master[67].sequencer;   
    sequencer.master_sequencer_D1868 =  pf_vf_mux_system_env_TB4_D3.master[68].sequencer;   
    sequencer.master_sequencer_D1869 =  pf_vf_mux_system_env_TB4_D3.master[69].sequencer;   
    sequencer.master_sequencer_D1870 =  pf_vf_mux_system_env_TB4_D3.master[70].sequencer;   
    sequencer.master_sequencer_D1871 =  pf_vf_mux_system_env_TB4_D3.master[71].sequencer;   
    sequencer.master_sequencer_D1872 =  pf_vf_mux_system_env_TB4_D3.master[72].sequencer;   
    sequencer.master_sequencer_D1873 =  pf_vf_mux_system_env_TB4_D3.master[73].sequencer;   
    sequencer.master_sequencer_D1874 =  pf_vf_mux_system_env_TB4_D3.master[74].sequencer;   
    sequencer.master_sequencer_D1875 =  pf_vf_mux_system_env_TB4_D3.master[75].sequencer;   
    sequencer.master_sequencer_D1876 =  pf_vf_mux_system_env_TB4_D3.master[76].sequencer;   
    sequencer.master_sequencer_D1877 =  pf_vf_mux_system_env_TB4_D3.master[77].sequencer;   
    sequencer.master_sequencer_D1878 =  pf_vf_mux_system_env_TB4_D3.master[78].sequencer;   
    sequencer.master_sequencer_D1879 =  pf_vf_mux_system_env_TB4_D3.master[79].sequencer;   
    sequencer.master_sequencer_D1880 =  pf_vf_mux_system_env_TB4_D3.master[80].sequencer;   
    sequencer.master_sequencer_D1881 =  pf_vf_mux_system_env_TB4_D3.master[81].sequencer;   
    sequencer.master_sequencer_D1882 =  pf_vf_mux_system_env_TB4_D3.master[82].sequencer;   
    sequencer.master_sequencer_D1883 =  pf_vf_mux_system_env_TB4_D3.master[83].sequencer;   
    sequencer.master_sequencer_D1884 =  pf_vf_mux_system_env_TB4_D3.master[84].sequencer;   
    sequencer.master_sequencer_D1885 =  pf_vf_mux_system_env_TB4_D3.master[85].sequencer;   
    sequencer.master_sequencer_D1886 =  pf_vf_mux_system_env_TB4_D3.master[86].sequencer;   
    sequencer.master_sequencer_D1887 =  pf_vf_mux_system_env_TB4_D3.master[87].sequencer;   
    sequencer.master_sequencer_D1888 =  pf_vf_mux_system_env_TB4_D3.master[88].sequencer;   
    sequencer.master_sequencer_D1889 =  pf_vf_mux_system_env_TB4_D3.master[89].sequencer;   
    sequencer.master_sequencer_D1890 =  pf_vf_mux_system_env_TB4_D3.master[90].sequencer;   
    sequencer.master_sequencer_D1891 =  pf_vf_mux_system_env_TB4_D3.master[91].sequencer;   
    sequencer.master_sequencer_D1892 =  pf_vf_mux_system_env_TB4_D3.master[92].sequencer;   
    sequencer.master_sequencer_D1893 =  pf_vf_mux_system_env_TB4_D3.master[93].sequencer;   
    sequencer.master_sequencer_D1894 =  pf_vf_mux_system_env_TB4_D3.master[94].sequencer;   
    sequencer.master_sequencer_D1895 =  pf_vf_mux_system_env_TB4_D3.master[95].sequencer;   
    sequencer.master_sequencer_D1896 =  pf_vf_mux_system_env_TB4_D3.master[96].sequencer;   
    sequencer.master_sequencer_D1897 =  pf_vf_mux_system_env_TB4_D3.master[97].sequencer;   
    sequencer.master_sequencer_D1898 =  pf_vf_mux_system_env_TB4_D3.master[98].sequencer;   
    sequencer.master_sequencer_D1899 =  pf_vf_mux_system_env_TB4_D3.master[99].sequencer;   
    sequencer.master_sequencer_D1900 =  pf_vf_mux_system_env_TB4_D3.master[100].sequencer;   
    sequencer.master_sequencer_D1901 =  pf_vf_mux_system_env_TB4_D3.master[101].sequencer;   
    sequencer.master_sequencer_D1902 =  pf_vf_mux_system_env_TB4_D3.master[102].sequencer;   
    sequencer.master_sequencer_D1903 =  pf_vf_mux_system_env_TB4_D3.master[103].sequencer;   
    sequencer.master_sequencer_D1904 =  pf_vf_mux_system_env_TB4_D3.master[104].sequencer;   
    sequencer.master_sequencer_D1905 =  pf_vf_mux_system_env_TB4_D3.master[105].sequencer;   
    sequencer.master_sequencer_D1906 =  pf_vf_mux_system_env_TB4_D3.master[106].sequencer;   
    sequencer.master_sequencer_D1907 =  pf_vf_mux_system_env_TB4_D3.master[107].sequencer;   
    sequencer.master_sequencer_D1908 =  pf_vf_mux_system_env_TB4_D3.master[108].sequencer;   
    sequencer.master_sequencer_D1909 =  pf_vf_mux_system_env_TB4_D3.master[109].sequencer;   
    sequencer.master_sequencer_D1910 =  pf_vf_mux_system_env_TB4_D3.master[110].sequencer;   
    sequencer.master_sequencer_D1911 =  pf_vf_mux_system_env_TB4_D3.master[111].sequencer;   
    sequencer.master_sequencer_D1912 =  pf_vf_mux_system_env_TB4_D3.master[112].sequencer;   
    sequencer.master_sequencer_D1913 =  pf_vf_mux_system_env_TB4_D3.master[113].sequencer;   
    sequencer.master_sequencer_D1914 =  pf_vf_mux_system_env_TB4_D3.master[114].sequencer;   
    sequencer.master_sequencer_D1915 =  pf_vf_mux_system_env_TB4_D3.master[115].sequencer;   
    sequencer.master_sequencer_D1916 =  pf_vf_mux_system_env_TB4_D3.master[116].sequencer;   
    sequencer.master_sequencer_D1917 =  pf_vf_mux_system_env_TB4_D3.master[117].sequencer;   
    sequencer.master_sequencer_D1918 =  pf_vf_mux_system_env_TB4_D3.master[118].sequencer;   
    sequencer.master_sequencer_D1919 =  pf_vf_mux_system_env_TB4_D3.master[119].sequencer;   
    sequencer.master_sequencer_D1920 =  pf_vf_mux_system_env_TB4_D3.master[120].sequencer;   
    sequencer.master_sequencer_D1921 =  pf_vf_mux_system_env_TB4_D3.master[121].sequencer;   
    sequencer.master_sequencer_D1922 =  pf_vf_mux_system_env_TB4_D3.master[122].sequencer;   
    sequencer.master_sequencer_D1923 =  pf_vf_mux_system_env_TB4_D3.master[123].sequencer;   
    sequencer.master_sequencer_D1924 =  pf_vf_mux_system_env_TB4_D3.master[124].sequencer;   
    sequencer.master_sequencer_D1925 =  pf_vf_mux_system_env_TB4_D3.master[125].sequencer;   
    sequencer.master_sequencer_D1926 =  pf_vf_mux_system_env_TB4_D3.master[126].sequencer;   
    sequencer.master_sequencer_D1927 =  pf_vf_mux_system_env_TB4_D3.master[127].sequencer;   
    sequencer.master_sequencer_D1928 =  pf_vf_mux_system_env_TB4_D3.master[128].sequencer;   
    sequencer.master_sequencer_D1929 =  pf_vf_mux_system_env_TB4_D3.master[129].sequencer;   
    sequencer.master_sequencer_D1930 =  pf_vf_mux_system_env_TB4_D3.master[130].sequencer;   
    sequencer.master_sequencer_D1931 =  pf_vf_mux_system_env_TB4_D3.master[131].sequencer;   
    sequencer.master_sequencer_D1932 =  pf_vf_mux_system_env_TB4_D3.master[132].sequencer;   
    sequencer.master_sequencer_D1933 =  pf_vf_mux_system_env_TB4_D3.master[133].sequencer;   
    sequencer.master_sequencer_D1934 =  pf_vf_mux_system_env_TB4_D3.master[134].sequencer;   
    sequencer.master_sequencer_D1935 =  pf_vf_mux_system_env_TB4_D3.master[135].sequencer;   
    sequencer.master_sequencer_D1936 =  pf_vf_mux_system_env_TB4_D3.master[136].sequencer;   
    sequencer.master_sequencer_D1937 =  pf_vf_mux_system_env_TB4_D3.master[137].sequencer;   
    sequencer.master_sequencer_D1938 =  pf_vf_mux_system_env_TB4_D3.master[138].sequencer;   
    sequencer.master_sequencer_D1939 =  pf_vf_mux_system_env_TB4_D3.master[139].sequencer;   
    sequencer.master_sequencer_D1940 =  pf_vf_mux_system_env_TB4_D3.master[140].sequencer;   
    sequencer.master_sequencer_D1941 =  pf_vf_mux_system_env_TB4_D3.master[141].sequencer;   
    sequencer.master_sequencer_D1942 =  pf_vf_mux_system_env_TB4_D3.master[142].sequencer;   
    sequencer.master_sequencer_D1943 =  pf_vf_mux_system_env_TB4_D3.master[143].sequencer;   
    sequencer.master_sequencer_D1944 =  pf_vf_mux_system_env_TB4_D3.master[144].sequencer;   
    sequencer.master_sequencer_D1945 =  pf_vf_mux_system_env_TB4_D3.master[145].sequencer;   
    sequencer.master_sequencer_D1946 =  pf_vf_mux_system_env_TB4_D3.master[146].sequencer;   
    sequencer.master_sequencer_D1947 =  pf_vf_mux_system_env_TB4_D3.master[147].sequencer;   
    sequencer.master_sequencer_D1948 =  pf_vf_mux_system_env_TB4_D3.master[148].sequencer;   
    sequencer.master_sequencer_D1949 =  pf_vf_mux_system_env_TB4_D3.master[149].sequencer;   
    sequencer.master_sequencer_D1950 =  pf_vf_mux_system_env_TB4_D3.master[150].sequencer;   
    sequencer.master_sequencer_D1951 =  pf_vf_mux_system_env_TB4_D3.master[151].sequencer;   
    sequencer.master_sequencer_D1952 =  pf_vf_mux_system_env_TB4_D3.master[152].sequencer;   
    sequencer.master_sequencer_D1953 =  pf_vf_mux_system_env_TB4_D3.master[153].sequencer;   
    sequencer.master_sequencer_D1954 =  pf_vf_mux_system_env_TB4_D3.master[154].sequencer;   
    sequencer.master_sequencer_D1955 =  pf_vf_mux_system_env_TB4_D3.master[155].sequencer;   
    sequencer.master_sequencer_D1956 =  pf_vf_mux_system_env_TB4_D3.master[156].sequencer;   
    sequencer.master_sequencer_D1957 =  pf_vf_mux_system_env_TB4_D3.master[157].sequencer;   
    sequencer.master_sequencer_D1958 =  pf_vf_mux_system_env_TB4_D3.master[158].sequencer;   
    sequencer.master_sequencer_D1959 =  pf_vf_mux_system_env_TB4_D3.master[159].sequencer;   
    sequencer.master_sequencer_D1960 =  pf_vf_mux_system_env_TB4_D3.master[160].sequencer;   
    sequencer.master_sequencer_D1961 =  pf_vf_mux_system_env_TB4_D3.master[161].sequencer;   
    sequencer.master_sequencer_D1962 =  pf_vf_mux_system_env_TB4_D3.master[162].sequencer;   
    sequencer.master_sequencer_D1963 =  pf_vf_mux_system_env_TB4_D3.master[163].sequencer;   
    sequencer.master_sequencer_D1964 =  pf_vf_mux_system_env_TB4_D3.master[164].sequencer;   
    sequencer.master_sequencer_D1965 =  pf_vf_mux_system_env_TB4_D3.master[165].sequencer;   
    sequencer.master_sequencer_D1966 =  pf_vf_mux_system_env_TB4_D3.master[166].sequencer;   
    sequencer.master_sequencer_D1967 =  pf_vf_mux_system_env_TB4_D3.master[167].sequencer;   
    sequencer.master_sequencer_D1968 =  pf_vf_mux_system_env_TB4_D3.master[168].sequencer;   
    sequencer.master_sequencer_D1969 =  pf_vf_mux_system_env_TB4_D3.master[169].sequencer;   
    sequencer.master_sequencer_D1970 =  pf_vf_mux_system_env_TB4_D3.master[170].sequencer;   
    sequencer.master_sequencer_D1971 =  pf_vf_mux_system_env_TB4_D3.master[171].sequencer;   
    sequencer.master_sequencer_D1972 =  pf_vf_mux_system_env_TB4_D3.master[172].sequencer;   
    sequencer.master_sequencer_D1973 =  pf_vf_mux_system_env_TB4_D3.master[173].sequencer;   
    sequencer.master_sequencer_D1974 =  pf_vf_mux_system_env_TB4_D3.master[174].sequencer;   
    sequencer.master_sequencer_D1975 =  pf_vf_mux_system_env_TB4_D3.master[175].sequencer;   
    sequencer.master_sequencer_D1976 =  pf_vf_mux_system_env_TB4_D3.master[176].sequencer;   
    sequencer.master_sequencer_D1977 =  pf_vf_mux_system_env_TB4_D3.master[177].sequencer;   
    sequencer.master_sequencer_D1978 =  pf_vf_mux_system_env_TB4_D3.master[178].sequencer;   
    sequencer.master_sequencer_D1979 =  pf_vf_mux_system_env_TB4_D3.master[179].sequencer;   
    sequencer.master_sequencer_D1980 =  pf_vf_mux_system_env_TB4_D3.master[180].sequencer;   
    sequencer.master_sequencer_D1981 =  pf_vf_mux_system_env_TB4_D3.master[181].sequencer;   
    sequencer.master_sequencer_D1982 =  pf_vf_mux_system_env_TB4_D3.master[182].sequencer;   
    sequencer.master_sequencer_D1983 =  pf_vf_mux_system_env_TB4_D3.master[183].sequencer;   
    sequencer.master_sequencer_D1984 =  pf_vf_mux_system_env_TB4_D3.master[184].sequencer;   
    sequencer.master_sequencer_D1985 =  pf_vf_mux_system_env_TB4_D3.master[185].sequencer;   
    sequencer.master_sequencer_D1986 =  pf_vf_mux_system_env_TB4_D3.master[186].sequencer;   
    sequencer.master_sequencer_D1987 =  pf_vf_mux_system_env_TB4_D3.master[187].sequencer;   
    sequencer.master_sequencer_D1988 =  pf_vf_mux_system_env_TB4_D3.master[188].sequencer;   
    sequencer.master_sequencer_D1989 =  pf_vf_mux_system_env_TB4_D3.master[189].sequencer;   
    sequencer.master_sequencer_D1990 =  pf_vf_mux_system_env_TB4_D3.master[190].sequencer;   
    sequencer.master_sequencer_D1991 =  pf_vf_mux_system_env_TB4_D3.master[191].sequencer;   
    sequencer.master_sequencer_D1992 =  pf_vf_mux_system_env_TB4_D3.master[192].sequencer;   
    sequencer.master_sequencer_D1993 =  pf_vf_mux_system_env_TB4_D3.master[193].sequencer;   
    sequencer.master_sequencer_D1994 =  pf_vf_mux_system_env_TB4_D3.master[194].sequencer;   
    sequencer.master_sequencer_D1995 =  pf_vf_mux_system_env_TB4_D3.master[195].sequencer;   
    sequencer.master_sequencer_D1996 =  pf_vf_mux_system_env_TB4_D3.master[196].sequencer;   
    sequencer.master_sequencer_D1997 =  pf_vf_mux_system_env_TB4_D3.master[197].sequencer;   
    sequencer.master_sequencer_D1998 =  pf_vf_mux_system_env_TB4_D3.master[198].sequencer;   
    sequencer.master_sequencer_D1999 =  pf_vf_mux_system_env_TB4_D3.master[199].sequencer;   
    sequencer.master_sequencer_D2000 =  pf_vf_mux_system_env_TB4_D3.master[200].sequencer;   
    sequencer.master_sequencer_D2001 =  pf_vf_mux_system_env_TB4_D3.master[201].sequencer;   
    sequencer.master_sequencer_D2002 =  pf_vf_mux_system_env_TB4_D3.master[202].sequencer;   
    sequencer.master_sequencer_D2003 =  pf_vf_mux_system_env_TB4_D3.master[203].sequencer;   
    sequencer.master_sequencer_D2004 =  pf_vf_mux_system_env_TB4_D3.master[204].sequencer;   
    sequencer.master_sequencer_D2005 =  pf_vf_mux_system_env_TB4_D3.master[205].sequencer;   
    sequencer.master_sequencer_D2006 =  pf_vf_mux_system_env_TB4_D3.master[206].sequencer;   
    sequencer.master_sequencer_D2007 =  pf_vf_mux_system_env_TB4_D3.master[207].sequencer;   
    sequencer.master_sequencer_D2008 =  pf_vf_mux_system_env_TB4_D3.master[208].sequencer;   
    sequencer.master_sequencer_D2009 =  pf_vf_mux_system_env_TB4_D3.master[209].sequencer;   
    sequencer.master_sequencer_D2010 =  pf_vf_mux_system_env_TB4_D3.master[210].sequencer;   
    sequencer.master_sequencer_D2011 =  pf_vf_mux_system_env_TB4_D3.master[211].sequencer;   
    sequencer.master_sequencer_D2012 =  pf_vf_mux_system_env_TB4_D3.master[212].sequencer;   
    sequencer.master_sequencer_D2013 =  pf_vf_mux_system_env_TB4_D3.master[213].sequencer;   
    sequencer.master_sequencer_D2014 =  pf_vf_mux_system_env_TB4_D3.master[214].sequencer;   
    sequencer.master_sequencer_D2015 =  pf_vf_mux_system_env_TB4_D3.master[215].sequencer;   
    sequencer.master_sequencer_D2016 =  pf_vf_mux_system_env_TB4_D3.master[216].sequencer;   
    sequencer.master_sequencer_D2017 =  pf_vf_mux_system_env_TB4_D3.master[217].sequencer;   
    sequencer.master_sequencer_D2018 =  pf_vf_mux_system_env_TB4_D3.master[218].sequencer;   
    sequencer.master_sequencer_D2019 =  pf_vf_mux_system_env_TB4_D3.master[219].sequencer;   
    sequencer.master_sequencer_D2020 =  pf_vf_mux_system_env_TB4_D3.master[220].sequencer;   
    sequencer.master_sequencer_D2021 =  pf_vf_mux_system_env_TB4_D3.master[221].sequencer;   
    sequencer.master_sequencer_D2022 =  pf_vf_mux_system_env_TB4_D3.master[222].sequencer;   
    sequencer.master_sequencer_D2023 =  pf_vf_mux_system_env_TB4_D3.master[223].sequencer;   
    sequencer.master_sequencer_D2024 =  pf_vf_mux_system_env_TB4_D3.master[224].sequencer;   
    sequencer.master_sequencer_D2025 =  pf_vf_mux_system_env_TB4_D3.master[225].sequencer;   
    sequencer.master_sequencer_D2026 =  pf_vf_mux_system_env_TB4_D3.master[226].sequencer;   
    sequencer.master_sequencer_D2027 =  pf_vf_mux_system_env_TB4_D3.master[227].sequencer;   
    sequencer.master_sequencer_D2028 =  pf_vf_mux_system_env_TB4_D3.master[228].sequencer;   
    sequencer.master_sequencer_D2029 =  pf_vf_mux_system_env_TB4_D3.master[229].sequencer;   
    sequencer.master_sequencer_D2030 =  pf_vf_mux_system_env_TB4_D3.master[230].sequencer;   
    sequencer.master_sequencer_D2031 =  pf_vf_mux_system_env_TB4_D3.master[231].sequencer;   
    sequencer.master_sequencer_D2032 =  pf_vf_mux_system_env_TB4_D3.master[232].sequencer;   
    sequencer.master_sequencer_D2033 =  pf_vf_mux_system_env_TB4_D3.master[233].sequencer;   
    sequencer.master_sequencer_D2034 =  pf_vf_mux_system_env_TB4_D3.master[234].sequencer;   
    sequencer.master_sequencer_D2035 =  pf_vf_mux_system_env_TB4_D3.master[235].sequencer;   
    sequencer.master_sequencer_D2036 =  pf_vf_mux_system_env_TB4_D3.master[236].sequencer;   
    sequencer.master_sequencer_D2037 =  pf_vf_mux_system_env_TB4_D3.master[237].sequencer;   
    sequencer.master_sequencer_D2038 =  pf_vf_mux_system_env_TB4_D3.master[238].sequencer;   
    sequencer.master_sequencer_D2039 =  pf_vf_mux_system_env_TB4_D3.master[239].sequencer;   
    sequencer.master_sequencer_D2040 =  pf_vf_mux_system_env_TB4_D3.master[240].sequencer;   
    sequencer.master_sequencer_D2041 =  pf_vf_mux_system_env_TB4_D3.master[241].sequencer;   
    sequencer.master_sequencer_D2042 =  pf_vf_mux_system_env_TB4_D3.master[242].sequencer;   
    sequencer.master_sequencer_D2043 =  pf_vf_mux_system_env_TB4_D3.master[243].sequencer;   
    sequencer.master_sequencer_D2044 =  pf_vf_mux_system_env_TB4_D3.master[244].sequencer;   
    sequencer.master_sequencer_D2045 =  pf_vf_mux_system_env_TB4_D3.master[245].sequencer;   
    sequencer.master_sequencer_D2046 =  pf_vf_mux_system_env_TB4_D3.master[246].sequencer;   
    sequencer.master_sequencer_D2047 =  pf_vf_mux_system_env_TB4_D3.master[247].sequencer;   


    `endif

    `uvm_info("connect_phase", "Exiting...", UVM_LOW)
  endfunction : connect_phase

  virtual task run_phase(uvm_phase phase);
     super.run_phase(phase);
    `uvm_info("run_phase", "Exiting...", UVM_LOW)
  endtask : run_phase

 function AXIS_HOST_CFG();
      cfg_H.num_masters = 1;
      cfg_H.num_slaves  = 1 ;

      cfg_H.create_sub_cfgs(1,1);

      cfg_H.master_cfg[0].axi_interface_type = svt_axi_port_configuration::AXI4_STREAM;
      cfg_H.slave_cfg[0].axi_interface_type = svt_axi_port_configuration::AXI4_STREAM;

      cfg_H.master_cfg[0].tdata_width = 512;
      cfg_H.master_cfg[0].tuser_width = 10;
      cfg_H.master_cfg[0].is_active = 1;
      cfg_H.master_cfg[0].default_tready=1;
      cfg_H.master_cfg[0].tstrb_enable=0;
      cfg_H.master_cfg[0].tid_enable=0;
      cfg_H.master_cfg[0].tdest_enable=0;
      cfg_H.master_cfg[0].tlast_enable=1;

      cfg_H.slave_cfg[0].tdata_width = 512;
      cfg_H.slave_cfg[0].tuser_width = 10;
      cfg_H.slave_cfg[0].is_active = 0;
      cfg_H.slave_cfg[0].default_tready=1;
      cfg_H.slave_cfg[0].tstrb_enable=0;
      cfg_H.slave_cfg[0].tid_enable=0;
      cfg_H.slave_cfg[0].tdest_enable=0;
      cfg_H.slave_cfg[0].tlast_enable=1;
     `ifdef INVALID_PF_VF
      cfg_H.tready_watchdog_timeout=0;   // DUT is responding differently for different pf-vf-vf_active combinations, causing PASS/FAIL(Assertion)
     `endif
 endfunction
    
  function AXIS_DEVICE_CFG();
      `ifdef TB_CONFIG_4
	      int no_of_devices = 450;
      `else
	      int no_of_devices = 16;
      `endif
      cfg_D.num_masters = no_of_devices ;
      cfg_D.num_slaves  = no_of_devices ;
      cfg_D.create_sub_cfgs(no_of_devices,no_of_devices);
	    for(int i=0;i<no_of_devices;i++) begin
      cfg_D.master_cfg[i].axi_interface_type = svt_axi_port_configuration::AXI4_STREAM;
      cfg_D.slave_cfg[i].axi_interface_type = svt_axi_port_configuration::AXI4_STREAM;
      cfg_D.master_cfg[i].tdata_width = 512;
      cfg_D.master_cfg[i].tuser_width = 10;
      cfg_D.master_cfg[i].is_active = 1;
      cfg_D.master_cfg[i].default_tready=1;
      cfg_D.master_cfg[i].tstrb_enable=0;
      cfg_D.master_cfg[i].tid_enable=0;
      cfg_D.master_cfg[i].tdest_enable=0;
      cfg_D.master_cfg[i].tlast_enable=1;
      cfg_D.slave_cfg[i].tdata_width = 512;
      cfg_D.slave_cfg[i].tuser_width = 10;
      cfg_D.slave_cfg[i].is_active = 0;
      cfg_D.slave_cfg[i].default_tready=1;
      cfg_D.slave_cfg[i].tstrb_enable=0;
      cfg_D.slave_cfg[i].tid_enable=0;
      cfg_D.slave_cfg[i].tdest_enable=0;
      cfg_D.slave_cfg[i].tlast_enable=1;
      end
  endfunction

`ifndef TB_CONFIG_4
 `ifndef TB_CONFIG_1
   function AXIS_DEVICE_CFG_N();
       int no_of_devices ;
      `ifdef TB_CONFIG_2
         no_of_devices = 8;
      `elsif TB_CONFIG_3
         no_of_devices = 16;
      `endif
      cfg_DN.num_masters = no_of_devices ;
      cfg_DN.num_slaves  = no_of_devices ;
      cfg_DN.create_sub_cfgs(no_of_devices,no_of_devices);
	    for(int i=0;i<no_of_devices;i++) begin
      cfg_DN.master_cfg[i].axi_interface_type = svt_axi_port_configuration::AXI4_STREAM;
      cfg_DN.slave_cfg[i].axi_interface_type = svt_axi_port_configuration::AXI4_STREAM;
      cfg_DN.master_cfg[i].tdata_width = 512;
      cfg_DN.master_cfg[i].tuser_width = 10;
      cfg_DN.master_cfg[i].is_active = 1;
      cfg_DN.master_cfg[i].default_tready=1;
      cfg_DN.master_cfg[i].tstrb_enable=0;
      cfg_DN.master_cfg[i].tid_enable=0;
      cfg_DN.master_cfg[i].tdest_enable=0;
      cfg_DN.master_cfg[i].tlast_enable=1;
      cfg_DN.slave_cfg[i].tdata_width = 512;
      cfg_DN.slave_cfg[i].tuser_width = 10;
      cfg_DN.slave_cfg[i].is_active = 0;
      cfg_DN.slave_cfg[i].default_tready=1;
      cfg_DN.slave_cfg[i].tstrb_enable=0;
      cfg_DN.slave_cfg[i].tid_enable=0;
      cfg_DN.slave_cfg[i].tdest_enable=0;
      cfg_DN.slave_cfg[i].tlast_enable=1;
      end
  endfunction
 `endif  
`endif

`ifdef TB_CONFIG_4
  function AXIS_DEVICE_TB4_CFG();
	    int no_of_devices = 450;
      cfg_TB4_D0.num_masters = no_of_devices ;
      cfg_TB4_D0.num_slaves  = no_of_devices ;
      cfg_TB4_D0.create_sub_cfgs(no_of_devices,no_of_devices);
	    for(int i=0;i<no_of_devices;i++) begin
      cfg_TB4_D0.master_cfg[i].axi_interface_type = svt_axi_port_configuration::AXI4_STREAM;
      cfg_TB4_D0.slave_cfg[i].axi_interface_type = svt_axi_port_configuration::AXI4_STREAM;
      cfg_TB4_D0.master_cfg[i].tdata_width = 512;
      cfg_TB4_D0.master_cfg[i].tuser_width = 10;
      cfg_TB4_D0.master_cfg[i].is_active = 1;
      cfg_TB4_D0.master_cfg[i].default_tready=1;
      cfg_TB4_D0.master_cfg[i].tstrb_enable=0;
      cfg_TB4_D0.master_cfg[i].tid_enable=0;
      cfg_TB4_D0.master_cfg[i].tdest_enable=0;
      cfg_TB4_D0.master_cfg[i].tlast_enable=1;
      cfg_TB4_D0.slave_cfg[i].tdata_width = 512;
      cfg_TB4_D0.slave_cfg[i].tuser_width = 10;
      cfg_TB4_D0.slave_cfg[i].is_active = 0;
      cfg_TB4_D0.slave_cfg[i].default_tready=1;
      cfg_TB4_D0.slave_cfg[i].tstrb_enable=0;
      cfg_TB4_D0.slave_cfg[i].tid_enable=0;
      cfg_TB4_D0.slave_cfg[i].tdest_enable=0;
      cfg_TB4_D0.slave_cfg[i].tlast_enable=1;
			end
			cfg_TB4_D1.num_masters = no_of_devices ;
      cfg_TB4_D1.num_slaves  = no_of_devices ;
      cfg_TB4_D1.create_sub_cfgs(no_of_devices,no_of_devices);
	    for(int i=0;i<no_of_devices;i++) begin
      cfg_TB4_D1.master_cfg[i].axi_interface_type = svt_axi_port_configuration::AXI4_STREAM;
      cfg_TB4_D1.slave_cfg[i].axi_interface_type = svt_axi_port_configuration::AXI4_STREAM;
      cfg_TB4_D1.master_cfg[i].tdata_width = 512;
      cfg_TB4_D1.master_cfg[i].tuser_width = 10;
      cfg_TB4_D1.master_cfg[i].is_active = 1;
      cfg_TB4_D1.master_cfg[i].default_tready=1;
      cfg_TB4_D1.master_cfg[i].tstrb_enable=0;
      cfg_TB4_D1.master_cfg[i].tid_enable=0;
      cfg_TB4_D1.master_cfg[i].tdest_enable=0;
      cfg_TB4_D1.master_cfg[i].tlast_enable=1;
      cfg_TB4_D1.slave_cfg[i].tdata_width = 512;
      cfg_TB4_D1.slave_cfg[i].tuser_width = 10;
      cfg_TB4_D1.slave_cfg[i].is_active = 0;
      cfg_TB4_D1.slave_cfg[i].default_tready=1;
      cfg_TB4_D1.slave_cfg[i].tstrb_enable=0;
      cfg_TB4_D1.slave_cfg[i].tid_enable=0;
      cfg_TB4_D1.slave_cfg[i].tdest_enable=0;
      cfg_TB4_D1.slave_cfg[i].tlast_enable=1;
			end
			cfg_TB4_D2.num_masters = no_of_devices ;
      cfg_TB4_D2.num_slaves  = no_of_devices ;
      cfg_TB4_D2.create_sub_cfgs(no_of_devices,no_of_devices);
	    for(int i=0;i<no_of_devices;i++) begin
      cfg_TB4_D2.master_cfg[i].axi_interface_type = svt_axi_port_configuration::AXI4_STREAM;
      cfg_TB4_D2.slave_cfg[i].axi_interface_type = svt_axi_port_configuration::AXI4_STREAM;
      cfg_TB4_D2.master_cfg[i].tdata_width = 512;
      cfg_TB4_D2.master_cfg[i].tuser_width = 10;
      cfg_TB4_D2.master_cfg[i].is_active = 1;
      cfg_TB4_D2.master_cfg[i].default_tready=1;
      cfg_TB4_D2.master_cfg[i].tstrb_enable=0;
      cfg_TB4_D2.master_cfg[i].tid_enable=0;
      cfg_TB4_D2.master_cfg[i].tdest_enable=0;
      cfg_TB4_D2.master_cfg[i].tlast_enable=1;
      cfg_TB4_D2.slave_cfg[i].tdata_width = 512;
      cfg_TB4_D2.slave_cfg[i].tuser_width = 10;
      cfg_TB4_D2.slave_cfg[i].is_active = 0;
      cfg_TB4_D2.slave_cfg[i].default_tready=1;
      cfg_TB4_D2.slave_cfg[i].tstrb_enable=0;
      cfg_TB4_D2.slave_cfg[i].tid_enable=0;
      cfg_TB4_D2.slave_cfg[i].tdest_enable=0;
      cfg_TB4_D2.slave_cfg[i].tlast_enable=1;
			end
			cfg_TB4_D3.num_masters = no_of_devices ;
      cfg_TB4_D3.num_slaves  = no_of_devices ;
      cfg_TB4_D3.create_sub_cfgs(no_of_devices,no_of_devices);
	    for(int i=0;i<no_of_devices;i++) begin
      cfg_TB4_D3.master_cfg[i].axi_interface_type = svt_axi_port_configuration::AXI4_STREAM;
      cfg_TB4_D3.slave_cfg[i].axi_interface_type = svt_axi_port_configuration::AXI4_STREAM;
      cfg_TB4_D3.master_cfg[i].tdata_width = 512;
      cfg_TB4_D3.master_cfg[i].tuser_width = 10;
      cfg_TB4_D3.master_cfg[i].is_active = 1;
      cfg_TB4_D3.master_cfg[i].default_tready=1;
      cfg_TB4_D3.master_cfg[i].tstrb_enable=0;
      cfg_TB4_D3.master_cfg[i].tid_enable=0;
      cfg_TB4_D3.master_cfg[i].tdest_enable=0;
      cfg_TB4_D3.master_cfg[i].tlast_enable=1;
      cfg_TB4_D3.slave_cfg[i].tdata_width = 512;
      cfg_TB4_D3.slave_cfg[i].tuser_width = 10;
      cfg_TB4_D3.slave_cfg[i].is_active = 0;
      cfg_TB4_D3.slave_cfg[i].default_tready=1;
      cfg_TB4_D3.slave_cfg[i].tstrb_enable=0;
      cfg_TB4_D3.slave_cfg[i].tid_enable=0;
      cfg_TB4_D3.slave_cfg[i].tdest_enable=0;
      cfg_TB4_D3.slave_cfg[i].tlast_enable=1;
      end
  endfunction
`endif  

  
endclass

`endif // GUARD_pf_vf_mux_basic_env_SV
