// Copyright (C) 2023 Intel Corporation
// SPDX-License-Identifier: MIT

`define payload_generate(PF,VF,VA) \
          local_vf_active = ``VA``;\
          local_pf_num    = ``PF``;\
          local_vf_num    = ``VF``;\
          local_tlp_length = $urandom_range(1,64) ;\
          local_payload = 'h0;\
          local_my_payload = 'h0;\
          assert(std::randomize(random_value));\      
          for(int j=0; j < (local_tlp_length*32); j++) local_my_payload[j] = 1'b1;\
          local_payload = (random_value) & local_my_payload;\
          `uvm_info("body", $sformatf("TLP Length = %h and Payload = %h and Random Value generated = %h No of Trans = %d",local_tlp_length,local_payload,random_value,no_of_transactions),UVM_LOW)\
     
class pf_vf_mux_slave_fifo_error_seq extends uvm_sequence;
    
     rand bit local_vf_active       ;
     rand bit [2:0] local_pf_num    ;
     rand bit [10:0] local_vf_num   ;
     bit [9:0] local_tlp_length;
     bit [255:0] local_payload , random_value, local_my_payload;
     rand int no_of_transactions ;
     int num = 0;
    `uvm_object_utils(pf_vf_mux_slave_fifo_error_seq);

  /** Declare a typed sequencer object that the sequence can access */
  `uvm_declare_p_sequencer(pf_vf_mux_virtual_sequencer)


    function new (string name = "pf_vf_mux_slave_fifo_error_seq");
        super.new(name);
    endfunction : new

     virtual function void build_phase(uvm_phase phase);
        `uvm_info ("build_phase", "Entered PF Traffic Sequence Build Phase...",UVM_LOW);
      endfunction: build_phase


    task body();
        pf_vf_mux_request_sequence master_seq;
        super.body(); 
      	`uvm_info(get_name(), "Entering PF0 Traffic sequence...", UVM_LOW)
        `uvm_info(get_name(), "Starting master sequence on Device master sequencer", UVM_LOW)

     for(int i=0; i<no_of_transactions; i++)     
     begin//{    
     if (i==0)
       begin
       `uvm_info("body", "UNDERFLOW_FIFO_ERR_``PORT``", UVM_LOW) 
       force top_tb.pf_vf_mux_a.switch.M_mux[0].out_q.fifo_ren = 1;      //to check fifo_err for the case read after fifo_empty
       end 
     else force top_tb.pf_vf_mux_a.switch.M_mux[0].out_q.fifo_ren = 0;       
 
     if(top_tb.pf_vf_mux_a.switch.M_mux[0].out_q.full==1) begin          //to check fifo_err for the case write after fifo_full
         `uvm_info(get_name(), "Fifo full...", UVM_LOW)
         `uvm_info("body", "OVERFLOW_FIFO_ERR_``PORT``", UVM_LOW)
          force top_tb.pf_vf_mux_a.switch.M_mux[0].out_q.fifo_w = 1;
          @(posedge top_tb.pf_vf_mux_a.switch.M_mux[0].out_q.clk);
          force top_tb.pf_vf_mux_a.switch.M_mux[0].out_q.fifo_w = 0;
     end           
     else if (top_tb.pf_vf_mux_a.switch.M_mux[0].out_q.full==0)
	   `uvm_info(get_name(), "Fifo not full...", UVM_LOW)

     fork//{
         begin
           if(i<=(no_of_transactions/3)) 
             force top_tb.mx2ho_tx_remap.tready         =  1;
           else if ((i>=(no_of_transactions/3)) && (i<=(2*no_of_transactions/3)))
             force top_tb.mx2ho_tx_remap.tready         =  0; 
           else  
             force top_tb.mx2ho_tx_remap.tready         =  1; 
         end
        `ifndef TB_CONFIG_4 
         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'h0,'h0);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D0, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                      
                                                                                              })
           

            
         end
     
         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h1,'h0,'h0);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                      
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h2,'h0,'h0);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                      
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h3,'h0,'h0);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D3, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                     
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h4,'h0,'h0);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D4, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                     
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h5,'h0,'h0);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D5, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                     
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h6,'h0,'h0);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D6, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                      
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h7,'h0,'h0);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D7, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                      
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h0,'h0,'h1);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D8, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                    
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h1,'h0,'h1);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D9, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h2,'h0,'h1);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D10, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                     
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h3,'h0,'h1);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D11, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                    
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h4,'h0,'h1);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D12, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                   
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h5,'h0,'h1);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D13, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                      
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h6,'h0,'h1);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D14, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                      
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h7,'h0,'h1);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D15, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                      
                                                                                              })
           

         end
         `ifndef TB_CONFIG_1
         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h0,'h7FF,'h1);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D0, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                         direction   == 1'b1              ;
                                                                                      
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h1,'h7FF,'h1);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                      
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h2,'h7FF,'h1);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                      
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h3,'h7FF,'h1);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D3, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                      
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h4,'h7FF,'h1);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D4, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                      
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h5,'h7FF,'h1);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D5, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                      
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h6,'h7FF,'h1);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D6, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                      
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h7,'h7FF,'h1);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D7, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                      
                                                                                              })
           

         end
         `endif
     
         `ifdef TB_CONFIG_3
         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h0,`RANDOM_VF,'h1);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D8, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                      
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h1,`RANDOM_VF,'h1);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D9, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                      
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h2,`RANDOM_VF,'h1);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D10, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                      
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h3,`RANDOM_VF,'h1);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D11, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                      
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h4,`RANDOM_VF,'h1);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D12, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                      
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h5,`RANDOM_VF,'h1);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D13, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                      
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h6,`RANDOM_VF,'h1);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D14, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                      
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h7,`RANDOM_VF,'h1);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D15, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                      
                                                                                              })
           

         end
         `endif
       `endif

       `ifdef TB_CONFIG_4
        begin
        `payload_generate('h0,0,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D0, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,2,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,3,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D3, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,4,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D4, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,5,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D5, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,6,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D6, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,7,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D7, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,8,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D8, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,9,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D9, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,10,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D10, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,11,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D11, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,12,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D12, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,13,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D13, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,14,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D14, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,15,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D15, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,16,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D16, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,17,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D17, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,18,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D18, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,19,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D19, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,20,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D20, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,21,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D21, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,22,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D22, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,23,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D23, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,24,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D24, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,25,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D25, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,26,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D26, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,27,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D27, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,28,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D28, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,29,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D29, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,30,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D30, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,31,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D31, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,32,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D32, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,33,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D33, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,34,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D34, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,35,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D35, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,36,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D36, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,37,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D37, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,38,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D38, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,39,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D39, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,40,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D40, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,41,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D41, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,42,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D42, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,43,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D43, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,44,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D44, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,45,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D45, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,46,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D46, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,47,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D47, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,48,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D48, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,49,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D49, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,50,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D50, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,51,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D51, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,52,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D52, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,53,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D53, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,54,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D54, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,55,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D55, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,56,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D56, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,57,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D57, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,58,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D58, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,59,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D59, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,60,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D60, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,61,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D61, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,62,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D62, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,63,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D63, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,64,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D64, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,65,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D65, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,66,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D66, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,67,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D67, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,68,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D68, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,69,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D69, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,70,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D70, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,71,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D71, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,72,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D72, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,73,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D73, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,74,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D74, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,75,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D75, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,76,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D76, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,77,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D77, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,78,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D78, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,79,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D79, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,80,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D80, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,81,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D81, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,82,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D82, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,83,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D83, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,84,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D84, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,85,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D85, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,86,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D86, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,87,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D87, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,88,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D88, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,89,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D89, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,90,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D90, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,91,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D91, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,92,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D92, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,93,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D93, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,94,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D94, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,95,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D95, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,96,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D96, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,97,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D97, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,98,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D98, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,99,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D99, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,100,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D100, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,101,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D101, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,102,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D102, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,103,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D103, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,104,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D104, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,105,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D105, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,106,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D106, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,107,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D107, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,108,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D108, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,109,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D109, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,110,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D110, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,111,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D111, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,112,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D112, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,113,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D113, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,114,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D114, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,115,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D115, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,116,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D116, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,117,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D117, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,118,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D118, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,119,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D119, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,120,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D120, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,121,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D121, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,122,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D122, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,123,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D123, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,124,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D124, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,125,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D125, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,126,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D126, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,127,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D127, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,128,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D128, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,129,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D129, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,130,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D130, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,131,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D131, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,132,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D132, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,133,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D133, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,134,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D134, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,135,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D135, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,136,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D136, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,137,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D137, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,138,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D138, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,139,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D139, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,140,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D140, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,141,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D141, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,142,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D142, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,143,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D143, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,144,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D144, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,145,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D145, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,146,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D146, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,147,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D147, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,148,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D148, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,149,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D149, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,150,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D150, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,151,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D151, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,152,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D152, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,153,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D153, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,154,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D154, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,155,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D155, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,156,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D156, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,157,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D157, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,158,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D158, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,159,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D159, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,160,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D160, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,161,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D161, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,162,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D162, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,163,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D163, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,164,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D164, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,165,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D165, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,166,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D166, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,167,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D167, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,168,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D168, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,169,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D169, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,170,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D170, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,171,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D171, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,172,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D172, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,173,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D173, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,174,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D174, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,175,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D175, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,176,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D176, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,177,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D177, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,178,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D178, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,179,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D179, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,180,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D180, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,181,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D181, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,182,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D182, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,183,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D183, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,184,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D184, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,185,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D185, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,186,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D186, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,187,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D187, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,188,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D188, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,189,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D189, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,190,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D190, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,191,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D191, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,192,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D192, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,193,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D193, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,194,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D194, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,195,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D195, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,196,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D196, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,197,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D197, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,198,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D198, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,199,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D199, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,200,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D200, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,201,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D201, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,202,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D202, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,203,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D203, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,204,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D204, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,205,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D205, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,206,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D206, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,207,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D207, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,208,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D208, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,209,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D209, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,210,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D210, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,211,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D211, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,212,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D212, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,213,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D213, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,214,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D214, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,215,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D215, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,216,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D216, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,217,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D217, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,218,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D218, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,219,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D219, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,220,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D220, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,221,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D221, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,222,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D222, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,223,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D223, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,224,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D224, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,225,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D225, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,226,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D226, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,227,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D227, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,228,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D228, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,229,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D229, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,230,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D230, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,231,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D231, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,232,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D232, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,233,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D233, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,234,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D234, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,235,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D235, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,236,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D236, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,237,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D237, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,238,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D238, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,239,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D239, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,240,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D240, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,241,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D241, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,242,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D242, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,243,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D243, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,244,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D244, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,245,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D245, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,246,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D246, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,247,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D247, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,248,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D248, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,249,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D249, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,250,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D250, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,251,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D251, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,252,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D252, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,253,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D253, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,254,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D254, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,255,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D255, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,256,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D256, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,257,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D257, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,258,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D258, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,259,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D259, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,260,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D260, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,261,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D261, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,262,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D262, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,263,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D263, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,264,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D264, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,265,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D265, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,266,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D266, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,267,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D267, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,268,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D268, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,269,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D269, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,270,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D270, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,271,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D271, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,272,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D272, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,273,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D273, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,274,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D274, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,275,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D275, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,276,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D276, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,277,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D277, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,278,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D278, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,279,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D279, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,280,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D280, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,281,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D281, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,282,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D282, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,283,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D283, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,284,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D284, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,285,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D285, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,286,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D286, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,287,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D287, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,288,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D288, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,289,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D289, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,290,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D290, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,291,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D291, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,292,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D292, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,293,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D293, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,294,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D294, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,295,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D295, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,296,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D296, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,297,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D297, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,298,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D298, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,299,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D299, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,300,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D300, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,301,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D301, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,302,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D302, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,303,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D303, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,304,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D304, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,305,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D305, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,306,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D306, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,307,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D307, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,308,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D308, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,309,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D309, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,310,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D310, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,311,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D311, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,312,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D312, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,313,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D313, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,314,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D314, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,315,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D315, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,316,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D316, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,317,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D317, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,318,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D318, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,319,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D319, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,320,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D320, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,321,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D321, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,322,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D322, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,323,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D323, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,324,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D324, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,325,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D325, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,326,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D326, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,327,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D327, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,328,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D328, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,329,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D329, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,330,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D330, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,331,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D331, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,332,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D332, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,333,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D333, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,334,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D334, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,335,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D335, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,336,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D336, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,337,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D337, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,338,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D338, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,339,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D339, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,340,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D340, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,341,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D341, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,342,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D342, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,343,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D343, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,344,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D344, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,345,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D345, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,346,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D346, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,347,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D347, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,348,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D348, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,349,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D349, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,350,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D350, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,351,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D351, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,352,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D352, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,353,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D353, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,354,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D354, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,355,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D355, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,356,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D356, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,357,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D357, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,358,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D358, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,359,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D359, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,360,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D360, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,361,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D361, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,362,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D362, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,363,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D363, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,364,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D364, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,365,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D365, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,366,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D366, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,367,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D367, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,368,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D368, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,369,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D369, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,370,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D370, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,371,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D371, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,372,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D372, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,373,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D373, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,374,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D374, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,375,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D375, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,376,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D376, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,377,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D377, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,378,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D378, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,379,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D379, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,380,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D380, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,381,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D381, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,382,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D382, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,383,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D383, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,384,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D384, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,385,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D385, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,386,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D386, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,387,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D387, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,388,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D388, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,389,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D389, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,390,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D390, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,391,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D391, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,392,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D392, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,393,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D393, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,394,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D394, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,395,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D395, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,396,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D396, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,397,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D397, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,398,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D398, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,399,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D399, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,400,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D400, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,401,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D401, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,402,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D402, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,403,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D403, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,404,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D404, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,405,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D405, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,406,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D406, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,407,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D407, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,408,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D408, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,409,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D409, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,410,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D410, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,411,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D411, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,412,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D412, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,413,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D413, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,414,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D414, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,415,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D415, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,416,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D416, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,417,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D417, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,418,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D418, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,419,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D419, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,420,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D420, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,421,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D421, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,422,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D422, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,423,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D423, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,424,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D424, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,425,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D425, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,426,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D426, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,427,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D427, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,428,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D428, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,429,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D429, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,430,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D430, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,431,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D431, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,432,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D432, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,433,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D433, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,434,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D434, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,435,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D435, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,436,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D436, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,437,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D437, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,438,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D438, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,439,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D439, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,440,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D440, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,441,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D441, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,442,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D442, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,443,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D443, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,444,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D444, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,445,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D445, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,446,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D446, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,447,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D447, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,448,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D448, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,449,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D449, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,450,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D450, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,451,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D451, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,452,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D452, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,453,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D453, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,454,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D454, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,455,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D455, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,456,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D456, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,457,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D457, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,458,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D458, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,459,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D459, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,460,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D460, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,461,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D461, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,462,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D462, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,463,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D463, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,464,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D464, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,465,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D465, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,466,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D466, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,467,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D467, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,468,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D468, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,469,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D469, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,470,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D470, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,471,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D471, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,472,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D472, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,473,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D473, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,474,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D474, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,475,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D475, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,476,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D476, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,477,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D477, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,478,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D478, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,479,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D479, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,480,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D480, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,481,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D481, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,482,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D482, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,483,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D483, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,484,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D484, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,485,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D485, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,486,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D486, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,487,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D487, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,488,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D488, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,489,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D489, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,490,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D490, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,491,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D491, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,492,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D492, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,493,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D493, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,494,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D494, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,495,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D495, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,496,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D496, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,497,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D497, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,498,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D498, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,499,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D499, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,500,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D500, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,501,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D501, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,502,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D502, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,503,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D503, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,504,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D504, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,505,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D505, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,506,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D506, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,507,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D507, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,508,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D508, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,509,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D509, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,510,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D510, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,511,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D511, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,512,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D512, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,513,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D513, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,514,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D514, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,515,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D515, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,516,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D516, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,517,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D517, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,518,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D518, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,519,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D519, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,520,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D520, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,521,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D521, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,522,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D522, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,523,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D523, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,524,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D524, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,525,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D525, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,526,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D526, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,527,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D527, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,528,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D528, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,529,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D529, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,530,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D530, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,531,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D531, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,532,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D532, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,533,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D533, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,534,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D534, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,535,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D535, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,536,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D536, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,537,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D537, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,538,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D538, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,539,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D539, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,540,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D540, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,541,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D541, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,542,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D542, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,543,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D543, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,544,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D544, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,545,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D545, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,546,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D546, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,547,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D547, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,548,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D548, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,549,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D549, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,550,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D550, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,551,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D551, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,552,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D552, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,553,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D553, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,554,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D554, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,555,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D555, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,556,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D556, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,557,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D557, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,558,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D558, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,559,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D559, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,560,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D560, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,561,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D561, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,562,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D562, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,563,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D563, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,564,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D564, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,565,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D565, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,566,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D566, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,567,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D567, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,568,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D568, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,569,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D569, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,570,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D570, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,571,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D571, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,572,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D572, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,573,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D573, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,574,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D574, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,575,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D575, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,576,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D576, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,577,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D577, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,578,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D578, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,579,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D579, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,580,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D580, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,581,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D581, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,582,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D582, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,583,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D583, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,584,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D584, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,585,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D585, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,586,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D586, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,587,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D587, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,588,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D588, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,589,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D589, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,590,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D590, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,591,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D591, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,592,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D592, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,593,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D593, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,594,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D594, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,595,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D595, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,596,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D596, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,597,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D597, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,598,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D598, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,599,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D599, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,600,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D600, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,601,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D601, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,602,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D602, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,603,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D603, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,604,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D604, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,605,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D605, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,606,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D606, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,607,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D607, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,608,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D608, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,609,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D609, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,610,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D610, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,611,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D611, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,612,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D612, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,613,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D613, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,614,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D614, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,615,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D615, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,616,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D616, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,617,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D617, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,618,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D618, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,619,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D619, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,620,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D620, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,621,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D621, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,622,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D622, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,623,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D623, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,624,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D624, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,625,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D625, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,626,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D626, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,627,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D627, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,628,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D628, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,629,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D629, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,630,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D630, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,631,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D631, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,632,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D632, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,633,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D633, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,634,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D634, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,635,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D635, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,636,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D636, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,637,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D637, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,638,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D638, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,639,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D639, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,640,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D640, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,641,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D641, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,642,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D642, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,643,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D643, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,644,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D644, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,645,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D645, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,646,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D646, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,647,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D647, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,648,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D648, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,649,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D649, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,650,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D650, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,651,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D651, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,652,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D652, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,653,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D653, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,654,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D654, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,655,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D655, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,656,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D656, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,657,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D657, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,658,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D658, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,659,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D659, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,660,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D660, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,661,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D661, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,662,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D662, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,663,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D663, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,664,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D664, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,665,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D665, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,666,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D666, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,667,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D667, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,668,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D668, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,669,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D669, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,670,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D670, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,671,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D671, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,672,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D672, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,673,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D673, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,674,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D674, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,675,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D675, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,676,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D676, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,677,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D677, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,678,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D678, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,679,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D679, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,680,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D680, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,681,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D681, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,682,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D682, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,683,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D683, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,684,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D684, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,685,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D685, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,686,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D686, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,687,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D687, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,688,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D688, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,689,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D689, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,690,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D690, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,691,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D691, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,692,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D692, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,693,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D693, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,694,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D694, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,695,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D695, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,696,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D696, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,697,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D697, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,698,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D698, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,699,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D699, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,700,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D700, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,701,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D701, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,702,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D702, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,703,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D703, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,704,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D704, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,705,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D705, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,706,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D706, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,707,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D707, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,708,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D708, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,709,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D709, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,710,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D710, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,711,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D711, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,712,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D712, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,713,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D713, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,714,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D714, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,715,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D715, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,716,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D716, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,717,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D717, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,718,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D718, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,719,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D719, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,720,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D720, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,721,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D721, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,722,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D722, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,723,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D723, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,724,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D724, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,725,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D725, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,726,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D726, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,727,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D727, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,728,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D728, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,729,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D729, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,730,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D730, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,731,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D731, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,732,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D732, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,733,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D733, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,734,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D734, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,735,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D735, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,736,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D736, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,737,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D737, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,738,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D738, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,739,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D739, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,740,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D740, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,741,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D741, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,742,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D742, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,743,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D743, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,744,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D744, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,745,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D745, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,746,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D746, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,747,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D747, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,748,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D748, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,749,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D749, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,750,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D750, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,751,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D751, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,752,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D752, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,753,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D753, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,754,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D754, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,755,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D755, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,756,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D756, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,757,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D757, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,758,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D758, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,759,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D759, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,760,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D760, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,761,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D761, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,762,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D762, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,763,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D763, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,764,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D764, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,765,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D765, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,766,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D766, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,767,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D767, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,768,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D768, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,769,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D769, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,770,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D770, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,771,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D771, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,772,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D772, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,773,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D773, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,774,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D774, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,775,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D775, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,776,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D776, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,777,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D777, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,778,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D778, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,779,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D779, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,780,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D780, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,781,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D781, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,782,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D782, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,783,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D783, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,784,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D784, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,785,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D785, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,786,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D786, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,787,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D787, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,788,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D788, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,789,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D789, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,790,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D790, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,791,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D791, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,792,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D792, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,793,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D793, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,794,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D794, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,795,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D795, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,796,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D796, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,797,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D797, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,798,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D798, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,799,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D799, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,800,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D800, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,801,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D801, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,802,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D802, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,803,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D803, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,804,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D804, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,805,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D805, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,806,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D806, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,807,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D807, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,808,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D808, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,809,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D809, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,810,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D810, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,811,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D811, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,812,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D812, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,813,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D813, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,814,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D814, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,815,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D815, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,816,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D816, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,817,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D817, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,818,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D818, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,819,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D819, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,820,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D820, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,821,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D821, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,822,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D822, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,823,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D823, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,824,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D824, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,825,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D825, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,826,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D826, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,827,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D827, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,828,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D828, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,829,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D829, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,830,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D830, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,831,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D831, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,832,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D832, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,833,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D833, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,834,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D834, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,835,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D835, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,836,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D836, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,837,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D837, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,838,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D838, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,839,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D839, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,840,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D840, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,841,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D841, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,842,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D842, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,843,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D843, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,844,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D844, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,845,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D845, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,846,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D846, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,847,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D847, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,848,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D848, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,849,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D849, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,850,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D850, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,851,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D851, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,852,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D852, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,853,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D853, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,854,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D854, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,855,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D855, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,856,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D856, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,857,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D857, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,858,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D858, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,859,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D859, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,860,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D860, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,861,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D861, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,862,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D862, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,863,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D863, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,864,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D864, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,865,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D865, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,866,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D866, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,867,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D867, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,868,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D868, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,869,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D869, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,870,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D870, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,871,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D871, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,872,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D872, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,873,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D873, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,874,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D874, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,875,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D875, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,876,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D876, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,877,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D877, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,878,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D878, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,879,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D879, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,880,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D880, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,881,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D881, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,882,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D882, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,883,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D883, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,884,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D884, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,885,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D885, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,886,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D886, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,887,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D887, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,888,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D888, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,889,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D889, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,890,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D890, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,891,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D891, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,892,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D892, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,893,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D893, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,894,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D894, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,895,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D895, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,896,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D896, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,897,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D897, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,898,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D898, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,899,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D899, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,900,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D900, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,901,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D901, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,902,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D902, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,903,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D903, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,904,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D904, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,905,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D905, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,906,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D906, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,907,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D907, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,908,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D908, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,909,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D909, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,910,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D910, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,911,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D911, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,912,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D912, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,913,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D913, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,914,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D914, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,915,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D915, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,916,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D916, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,917,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D917, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,918,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D918, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,919,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D919, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,920,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D920, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,921,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D921, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,922,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D922, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,923,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D923, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,924,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D924, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,925,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D925, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,926,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D926, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,927,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D927, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,928,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D928, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,929,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D929, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,930,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D930, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,931,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D931, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,932,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D932, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,933,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D933, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,934,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D934, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,935,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D935, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,936,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D936, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,937,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D937, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,938,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D938, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,939,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D939, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,940,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D940, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,941,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D941, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,942,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D942, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,943,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D943, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,944,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D944, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,945,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D945, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,946,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D946, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,947,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D947, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,948,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D948, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,949,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D949, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,950,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D950, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,951,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D951, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,952,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D952, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,953,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D953, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,954,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D954, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,955,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D955, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,956,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D956, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,957,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D957, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,958,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D958, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,959,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D959, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,960,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D960, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,961,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D961, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,962,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D962, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,963,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D963, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,964,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D964, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,965,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D965, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,966,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D966, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,967,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D967, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,968,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D968, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,969,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D969, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,970,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D970, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,971,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D971, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,972,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D972, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,973,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D973, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,974,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D974, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,975,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D975, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,976,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D976, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,977,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D977, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,978,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D978, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,979,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D979, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,980,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D980, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,981,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D981, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,982,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D982, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,983,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D983, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,984,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D984, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,985,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D985, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,986,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D986, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,987,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D987, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,988,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D988, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,989,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D989, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,990,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D990, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,991,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D991, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,992,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D992, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,993,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D993, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,994,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D994, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,995,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D995, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,996,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D996, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,997,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D997, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,998,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D998, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,999,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D999, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1000,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1000, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1001,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1001, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1002,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1002, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1003,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1003, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1004,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1004, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1005,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1005, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1006,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1006, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1007,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1007, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1008,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1008, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1009,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1009, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1010,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1010, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1011,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1011, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1012,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1012, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1013,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1013, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1014,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1014, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1015,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1015, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1016,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1016, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1017,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1017, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1018,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1018, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1019,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1019, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1020,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1020, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1021,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1021, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1022,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1022, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1023,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1023, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1024,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1024, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1025,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1025, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1026,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1026, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1027,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1027, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1028,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1028, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1029,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1029, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1030,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1030, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1031,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1031, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1032,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1032, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1033,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1033, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1034,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1034, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1035,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1035, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1036,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1036, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1037,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1037, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1038,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1038, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1039,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1039, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1040,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1040, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1041,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1041, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1042,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1042, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1043,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1043, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1044,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1044, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1045,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1045, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1046,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1046, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1047,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1047, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1048,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1048, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1049,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1049, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1050,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1050, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1051,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1051, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1052,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1052, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1053,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1053, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1054,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1054, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1055,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1055, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1056,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1056, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1057,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1057, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1058,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1058, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1059,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1059, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1060,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1060, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1061,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1061, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1062,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1062, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1063,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1063, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1064,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1064, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1065,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1065, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1066,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1066, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1067,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1067, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1068,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1068, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1069,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1069, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1070,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1070, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1071,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1071, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1072,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1072, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1073,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1073, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1074,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1074, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1075,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1075, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1076,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1076, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1077,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1077, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1078,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1078, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1079,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1079, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1080,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1080, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1081,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1081, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1082,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1082, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1083,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1083, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1084,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1084, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1085,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1085, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1086,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1086, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1087,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1087, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1088,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1088, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1089,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1089, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1090,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1090, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1091,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1091, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1092,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1092, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1093,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1093, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1094,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1094, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1095,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1095, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1096,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1096, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1097,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1097, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1098,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1098, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1099,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1099, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1100,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1100, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1101,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1101, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1102,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1102, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1103,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1103, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1104,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1104, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1105,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1105, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1106,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1106, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1107,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1107, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1108,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1108, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1109,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1109, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1110,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1110, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1111,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1111, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1112,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1112, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1113,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1113, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1114,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1114, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1115,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1115, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1116,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1116, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1117,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1117, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1118,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1118, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1119,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1119, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1120,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1120, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1121,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1121, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1122,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1122, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1123,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1123, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1124,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1124, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1125,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1125, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1126,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1126, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1127,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1127, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1128,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1128, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1129,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1129, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1130,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1130, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1131,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1131, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1132,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1132, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1133,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1133, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1134,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1134, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1135,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1135, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1136,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1136, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1137,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1137, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1138,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1138, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1139,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1139, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1140,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1140, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1141,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1141, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1142,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1142, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1143,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1143, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1144,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1144, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1145,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1145, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1146,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1146, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1147,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1147, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1148,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1148, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1149,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1149, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1150,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1150, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1151,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1151, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1152,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1152, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1153,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1153, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1154,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1154, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1155,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1155, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1156,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1156, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1157,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1157, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1158,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1158, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1159,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1159, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1160,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1160, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1161,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1161, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1162,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1162, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1163,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1163, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1164,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1164, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1165,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1165, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1166,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1166, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1167,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1167, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1168,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1168, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1169,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1169, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1170,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1170, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1171,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1171, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1172,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1172, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1173,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1173, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1174,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1174, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1175,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1175, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1176,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1176, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1177,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1177, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1178,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1178, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1179,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1179, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1180,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1180, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1181,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1181, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1182,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1182, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1183,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1183, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1184,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1184, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1185,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1185, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1186,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1186, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1187,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1187, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1188,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1188, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1189,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1189, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1190,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1190, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1191,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1191, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1192,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1192, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1193,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1193, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1194,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1194, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1195,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1195, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1196,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1196, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1197,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1197, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1198,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1198, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1199,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1199, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1200,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1200, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1201,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1201, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1202,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1202, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1203,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1203, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1204,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1204, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1205,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1205, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1206,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1206, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1207,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1207, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1208,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1208, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1209,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1209, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1210,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1210, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1211,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1211, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1212,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1212, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1213,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1213, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1214,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1214, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1215,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1215, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1216,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1216, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1217,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1217, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1218,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1218, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1219,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1219, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1220,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1220, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1221,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1221, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1222,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1222, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1223,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1223, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1224,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1224, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1225,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1225, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1226,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1226, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1227,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1227, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1228,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1228, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1229,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1229, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1230,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1230, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1231,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1231, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1232,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1232, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1233,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1233, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1234,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1234, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1235,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1235, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1236,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1236, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1237,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1237, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1238,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1238, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1239,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1239, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1240,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1240, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1241,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1241, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1242,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1242, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1243,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1243, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1244,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1244, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1245,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1245, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1246,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1246, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1247,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1247, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1248,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1248, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1249,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1249, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1250,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1250, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1251,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1251, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1252,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1252, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1253,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1253, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1254,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1254, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1255,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1255, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1256,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1256, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1257,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1257, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1258,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1258, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1259,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1259, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1260,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1260, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1261,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1261, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1262,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1262, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1263,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1263, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1264,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1264, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1265,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1265, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1266,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1266, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1267,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1267, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1268,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1268, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1269,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1269, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1270,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1270, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1271,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1271, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1272,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1272, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1273,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1273, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1274,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1274, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1275,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1275, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1276,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1276, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1277,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1277, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1278,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1278, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1279,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1279, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1280,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1280, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1281,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1281, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1282,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1282, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1283,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1283, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1284,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1284, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1285,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1285, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1286,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1286, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1287,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1287, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1288,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1288, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1289,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1289, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1290,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1290, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1291,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1291, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1292,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1292, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1293,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1293, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1294,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1294, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1295,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1295, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1296,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1296, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1297,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1297, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1298,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1298, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1299,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1299, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1300,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1300, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1301,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1301, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1302,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1302, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1303,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1303, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1304,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1304, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1305,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1305, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1306,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1306, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1307,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1307, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1308,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1308, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1309,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1309, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1310,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1310, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1311,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1311, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1312,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1312, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1313,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1313, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1314,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1314, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1315,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1315, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1316,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1316, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1317,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1317, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1318,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1318, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1319,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1319, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1320,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1320, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1321,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1321, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1322,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1322, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1323,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1323, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1324,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1324, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1325,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1325, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1326,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1326, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1327,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1327, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1328,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1328, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1329,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1329, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1330,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1330, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1331,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1331, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1332,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1332, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1333,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1333, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1334,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1334, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1335,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1335, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1336,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1336, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1337,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1337, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1338,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1338, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1339,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1339, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1340,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1340, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1341,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1341, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1342,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1342, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1343,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1343, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1344,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1344, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1345,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1345, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1346,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1346, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1347,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1347, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1348,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1348, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1349,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1349, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1350,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1350, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1351,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1351, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1352,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1352, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1353,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1353, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1354,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1354, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1355,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1355, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1356,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1356, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1357,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1357, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1358,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1358, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1359,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1359, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1360,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1360, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1361,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1361, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1362,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1362, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1363,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1363, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1364,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1364, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1365,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1365, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1366,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1366, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1367,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1367, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1368,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1368, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1369,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1369, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1370,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1370, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1371,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1371, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1372,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1372, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1373,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1373, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1374,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1374, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1375,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1375, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1376,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1376, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1377,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1377, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1378,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1378, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1379,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1379, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1380,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1380, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1381,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1381, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1382,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1382, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1383,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1383, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1384,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1384, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1385,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1385, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1386,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1386, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1387,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1387, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1388,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1388, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1389,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1389, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1390,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1390, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1391,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1391, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1392,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1392, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1393,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1393, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1394,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1394, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1395,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1395, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1396,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1396, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1397,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1397, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1398,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1398, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1399,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1399, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1400,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1400, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1401,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1401, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1402,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1402, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1403,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1403, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1404,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1404, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1405,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1405, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1406,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1406, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1407,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1407, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1408,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1408, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1409,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1409, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1410,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1410, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1411,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1411, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1412,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1412, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1413,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1413, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1414,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1414, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1415,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1415, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1416,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1416, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1417,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1417, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1418,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1418, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1419,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1419, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1420,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1420, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1421,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1421, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1422,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1422, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1423,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1423, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1424,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1424, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1425,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1425, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1426,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1426, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1427,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1427, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1428,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1428, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1429,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1429, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1430,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1430, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1431,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1431, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1432,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1432, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1433,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1433, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1434,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1434, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1435,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1435, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1436,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1436, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1437,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1437, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1438,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1438, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1439,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1439, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1440,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1440, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1441,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1441, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1442,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1442, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1443,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1443, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1444,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1444, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1445,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1445, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1446,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1446, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1447,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1447, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1448,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1448, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1449,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1449, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1450,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1450, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1451,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1451, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1452,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1452, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1453,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1453, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1454,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1454, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1455,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1455, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1456,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1456, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1457,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1457, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1458,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1458, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1459,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1459, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1460,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1460, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1461,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1461, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1462,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1462, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1463,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1463, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1464,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1464, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1465,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1465, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1466,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1466, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1467,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1467, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1468,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1468, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1469,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1469, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1470,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1470, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1471,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1471, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1472,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1472, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1473,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1473, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1474,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1474, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1475,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1475, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1476,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1476, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1477,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1477, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1478,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1478, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1479,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1479, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1480,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1480, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1481,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1481, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1482,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1482, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1483,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1483, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1484,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1484, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1485,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1485, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1486,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1486, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1487,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1487, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1488,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1488, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1489,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1489, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1490,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1490, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1491,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1491, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1492,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1492, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1493,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1493, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1494,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1494, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1495,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1495, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1496,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1496, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1497,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1497, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1498,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1498, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1499,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1499, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1500,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1500, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1501,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1501, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1502,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1502, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1503,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1503, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1504,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1504, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1505,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1505, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1506,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1506, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1507,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1507, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1508,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1508, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1509,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1509, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1510,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1510, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1511,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1511, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1512,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1512, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1513,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1513, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1514,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1514, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1515,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1515, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1516,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1516, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1517,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1517, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1518,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1518, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1519,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1519, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1520,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1520, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1521,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1521, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1522,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1522, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1523,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1523, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1524,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1524, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1525,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1525, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1526,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1526, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1527,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1527, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1528,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1528, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1529,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1529, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1530,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1530, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1531,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1531, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1532,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1532, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1533,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1533, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1534,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1534, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1535,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1535, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1536,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1536, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1537,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1537, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1538,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1538, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1539,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1539, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1540,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1540, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1541,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1541, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1542,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1542, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1543,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1543, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1544,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1544, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1545,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1545, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1546,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1546, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1547,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1547, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1548,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1548, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1549,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1549, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1550,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1550, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1551,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1551, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1552,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1552, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1553,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1553, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1554,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1554, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1555,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1555, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1556,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1556, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1557,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1557, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1558,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1558, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1559,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1559, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1560,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1560, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1561,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1561, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1562,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1562, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1563,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1563, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1564,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1564, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1565,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1565, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1566,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1566, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1567,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1567, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1568,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1568, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1569,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1569, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1570,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1570, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1571,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1571, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1572,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1572, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1573,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1573, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1574,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1574, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1575,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1575, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1576,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1576, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1577,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1577, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1578,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1578, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1579,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1579, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1580,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1580, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1581,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1581, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1582,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1582, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1583,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1583, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1584,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1584, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1585,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1585, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1586,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1586, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1587,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1587, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1588,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1588, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1589,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1589, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1590,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1590, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1591,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1591, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1592,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1592, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1593,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1593, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1594,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1594, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1595,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1595, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1596,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1596, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1597,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1597, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1598,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1598, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1599,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1599, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1600,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1600, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1601,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1601, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1602,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1602, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1603,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1603, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1604,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1604, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1605,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1605, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1606,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1606, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1607,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1607, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1608,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1608, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1609,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1609, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1610,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1610, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1611,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1611, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1612,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1612, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1613,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1613, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1614,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1614, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1615,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1615, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1616,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1616, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1617,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1617, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1618,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1618, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1619,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1619, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1620,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1620, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1621,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1621, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1622,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1622, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1623,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1623, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1624,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1624, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1625,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1625, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1626,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1626, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1627,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1627, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1628,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1628, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1629,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1629, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1630,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1630, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1631,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1631, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1632,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1632, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1633,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1633, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1634,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1634, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1635,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1635, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1636,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1636, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1637,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1637, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1638,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1638, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1639,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1639, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1640,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1640, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1641,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1641, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1642,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1642, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1643,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1643, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1644,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1644, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1645,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1645, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1646,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1646, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1647,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1647, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1648,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1648, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1649,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1649, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1650,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1650, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1651,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1651, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1652,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1652, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1653,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1653, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1654,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1654, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1655,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1655, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1656,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1656, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1657,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1657, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1658,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1658, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1659,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1659, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1660,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1660, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1661,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1661, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1662,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1662, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1663,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1663, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1664,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1664, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1665,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1665, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1666,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1666, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1667,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1667, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1668,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1668, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1669,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1669, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1670,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1670, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1671,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1671, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1672,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1672, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1673,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1673, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1674,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1674, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1675,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1675, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1676,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1676, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1677,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1677, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1678,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1678, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1679,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1679, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1680,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1680, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1681,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1681, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1682,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1682, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1683,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1683, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1684,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1684, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1685,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1685, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1686,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1686, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1687,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1687, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1688,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1688, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1689,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1689, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1690,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1690, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1691,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1691, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1692,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1692, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1693,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1693, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1694,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1694, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1695,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1695, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1696,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1696, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1697,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1697, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1698,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1698, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1699,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1699, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1700,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1700, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1701,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1701, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1702,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1702, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1703,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1703, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1704,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1704, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1705,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1705, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1706,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1706, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1707,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1707, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1708,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1708, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1709,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1709, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1710,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1710, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1711,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1711, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1712,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1712, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1713,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1713, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1714,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1714, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1715,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1715, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1716,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1716, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1717,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1717, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1718,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1718, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1719,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1719, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1720,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1720, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1721,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1721, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1722,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1722, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1723,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1723, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1724,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1724, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1725,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1725, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1726,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1726, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1727,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1727, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1728,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1728, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1729,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1729, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1730,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1730, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1731,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1731, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1732,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1732, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1733,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1733, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1734,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1734, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1735,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1735, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1736,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1736, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1737,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1737, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1738,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1738, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1739,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1739, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1740,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1740, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1741,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1741, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1742,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1742, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1743,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1743, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1744,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1744, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1745,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1745, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1746,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1746, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1747,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1747, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1748,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1748, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1749,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1749, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1750,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1750, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1751,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1751, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1752,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1752, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1753,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1753, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1754,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1754, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1755,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1755, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1756,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1756, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1757,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1757, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1758,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1758, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1759,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1759, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1760,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1760, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1761,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1761, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1762,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1762, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1763,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1763, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1764,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1764, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1765,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1765, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1766,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1766, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1767,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1767, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1768,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1768, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1769,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1769, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1770,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1770, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1771,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1771, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1772,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1772, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1773,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1773, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1774,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1774, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1775,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1775, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1776,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1776, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1777,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1777, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1778,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1778, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1779,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1779, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1780,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1780, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1781,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1781, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1782,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1782, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1783,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1783, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1784,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1784, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1785,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1785, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1786,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1786, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1787,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1787, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1788,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1788, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1789,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1789, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1790,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1790, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1791,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1791, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1792,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1792, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1793,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1793, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1794,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1794, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1795,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1795, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1796,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1796, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1797,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1797, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1798,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1798, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1799,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1799, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1800,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1800, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1801,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1801, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1802,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1802, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1803,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1803, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1804,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1804, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1805,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1805, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1806,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1806, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1807,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1807, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1808,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1808, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1809,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1809, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1810,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1810, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1811,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1811, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1812,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1812, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1813,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1813, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1814,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1814, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1815,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1815, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1816,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1816, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1817,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1817, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1818,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1818, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1819,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1819, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1820,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1820, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1821,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1821, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1822,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1822, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1823,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1823, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1824,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1824, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1825,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1825, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1826,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1826, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1827,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1827, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1828,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1828, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1829,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1829, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1830,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1830, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1831,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1831, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1832,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1832, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1833,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1833, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1834,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1834, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1835,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1835, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1836,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1836, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1837,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1837, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1838,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1838, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1839,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1839, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1840,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1840, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1841,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1841, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1842,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1842, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1843,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1843, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1844,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1844, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1845,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1845, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1846,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1846, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1847,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1847, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1848,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1848, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1849,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1849, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1850,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1850, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1851,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1851, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1852,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1852, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1853,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1853, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1854,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1854, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1855,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1855, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1856,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1856, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1857,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1857, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1858,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1858, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1859,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1859, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1860,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1860, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1861,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1861, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1862,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1862, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1863,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1863, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1864,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1864, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1865,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1865, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1866,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1866, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1867,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1867, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1868,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1868, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1869,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1869, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1870,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1870, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1871,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1871, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1872,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1872, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1873,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1873, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1874,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1874, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1875,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1875, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1876,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1876, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1877,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1877, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1878,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1878, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1879,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1879, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1880,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1880, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1881,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1881, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1882,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1882, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1883,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1883, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1884,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1884, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1885,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1885, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1886,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1886, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1887,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1887, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1888,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1888, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1889,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1889, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1890,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1890, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1891,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1891, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1892,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1892, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1893,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1893, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1894,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1894, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1895,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1895, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1896,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1896, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1897,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1897, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1898,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1898, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1899,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1899, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1900,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1900, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1901,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1901, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1902,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1902, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1903,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1903, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1904,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1904, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1905,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1905, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1906,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1906, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1907,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1907, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1908,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1908, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1909,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1909, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1910,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1910, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1911,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1911, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1912,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1912, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1913,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1913, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1914,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1914, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1915,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1915, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1916,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1916, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1917,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1917, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1918,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1918, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1919,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1919, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1920,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1920, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1921,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1921, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1922,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1922, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1923,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1923, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1924,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1924, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1925,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1925, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1926,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1926, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1927,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1927, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1928,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1928, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1929,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1929, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1930,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1930, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1931,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1931, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1932,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1932, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1933,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1933, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1934,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1934, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1935,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1935, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1936,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1936, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1937,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1937, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1938,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1938, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1939,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1939, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1940,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1940, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1941,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1941, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1942,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1942, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1943,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1943, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1944,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1944, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1945,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1945, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1946,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1946, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1947,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1947, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1948,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1948, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1949,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1949, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1950,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1950, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1951,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1951, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1952,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1952, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1953,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1953, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1954,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1954, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1955,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1955, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1956,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1956, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1957,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1957, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1958,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1958, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1959,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1959, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1960,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1960, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1961,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1961, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1962,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1962, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1963,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1963, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1964,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1964, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1965,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1965, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1966,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1966, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1967,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1967, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1968,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1968, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1969,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1969, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1970,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1970, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1971,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1971, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1972,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1972, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1973,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1973, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1974,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1974, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1975,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1975, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1976,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1976, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1977,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1977, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1978,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1978, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1979,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1979, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1980,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1980, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1981,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1981, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1982,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1982, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1983,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1983, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1984,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1984, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1985,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1985, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1986,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1986, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1987,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1987, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1988,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1988, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1989,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1989, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1990,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1990, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1991,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1991, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1992,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1992, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1993,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1993, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1994,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1994, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1995,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1995, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1996,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1996, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1997,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1997, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1998,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1998, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,1999,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1999, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,2000,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2000, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,2001,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2001, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,2002,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2002, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,2003,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2003, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,2004,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2004, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,2005,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2005, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,2006,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2006, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,2007,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2007, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,2008,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2008, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,2009,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2009, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,2010,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2010, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,2011,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2011, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,2012,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2012, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,2013,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2013, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,2014,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2014, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,2015,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2015, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,2016,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2016, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,2017,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2017, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,2018,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2018, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,2019,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2019, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,2020,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2020, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,2021,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2021, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,2022,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2022, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,2023,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2023, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,2024,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2024, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,2025,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2025, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,2026,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2026, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,2027,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2027, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,2028,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2028, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,2029,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2029, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,2030,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2030, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,2031,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2031, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,2032,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2032, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,2033,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2033, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,2034,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2034, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,2035,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2035, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,2036,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2036, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,2037,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2037, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,2038,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2038, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,2039,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2039, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,2040,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2040, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,2041,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2041, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,2042,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2042, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,2043,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2043, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,2044,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2044, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,2045,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2045, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,2046,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2046, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end
        begin
        `payload_generate('h0,2047,'h1);
        `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2047, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        end

       `endif

join_none
wait fork;//}
end//}
    `uvm_info(get_name(), "Exiting sequence...", UVM_LOW)
    endtask : body

endclass
