// Copyright (C) 2023 Intel Corporation
// SPDX-License-Identifier: MIT

fork	

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d0,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D0, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d2,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d3,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D3, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d4,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D4, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d5,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D5, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d6,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D6, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d7,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D7, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d8,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D8, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d9,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D9, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d10,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D10, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d11,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D11, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d12,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D12, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d13,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D13, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d14,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D14, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d15,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D15, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d16,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D16, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d17,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D17, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d18,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D18, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d19,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D19, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d20,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D20, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d21,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D21, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d22,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D22, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d23,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D23, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d24,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D24, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d25,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D25, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d26,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D26, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d27,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D27, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d28,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D28, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d29,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D29, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d30,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D30, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d31,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D31, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d32,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D32, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d33,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D33, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d34,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D34, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d35,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D35, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d36,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D36, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d37,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D37, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d38,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D38, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d39,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D39, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d40,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D40, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d41,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D41, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d42,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D42, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d43,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D43, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d44,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D44, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d45,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D45, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d46,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D46, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d47,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D47, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d48,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D48, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d49,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D49, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d50,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D50, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d51,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D51, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d52,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D52, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d53,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D53, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d54,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D54, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d55,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D55, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d56,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D56, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d57,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D57, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d58,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D58, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d59,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D59, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d60,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D60, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d61,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D61, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d62,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D62, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d63,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D63, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d64,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D64, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d65,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D65, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d66,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D66, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d67,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D67, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d68,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D68, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d69,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D69, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d70,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D70, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d71,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D71, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d72,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D72, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d73,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D73, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d74,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D74, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d75,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D75, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d76,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D76, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d77,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D77, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d78,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D78, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d79,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D79, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d80,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D80, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d81,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D81, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d82,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D82, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d83,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D83, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d84,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D84, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d85,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D85, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d86,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D86, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d87,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D87, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d88,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D88, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d89,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D89, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d90,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D90, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d91,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D91, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d92,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D92, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d93,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D93, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d94,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D94, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d95,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D95, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d96,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D96, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d97,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D97, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d98,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D98, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d99,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D99, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d100,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D100, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d101,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D101, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d102,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D102, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d103,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D103, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d104,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D104, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d105,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D105, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d106,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D106, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d107,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D107, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d108,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D108, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d109,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D109, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d110,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D110, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d111,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D111, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d112,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D112, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d113,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D113, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d114,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D114, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d115,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D115, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d116,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D116, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d117,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D117, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d118,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D118, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d119,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D119, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d120,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D120, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d121,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D121, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d122,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D122, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d123,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D123, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d124,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D124, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d125,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D125, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d126,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D126, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d127,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D127, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d128,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D128, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d129,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D129, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d130,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D130, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d131,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D131, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d132,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D132, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d133,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D133, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d134,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D134, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d135,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D135, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d136,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D136, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d137,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D137, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d138,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D138, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d139,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D139, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d140,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D140, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d141,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D141, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d142,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D142, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d143,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D143, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d144,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D144, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d145,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D145, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d146,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D146, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d147,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D147, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d148,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D148, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d149,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D149, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d150,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D150, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d151,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D151, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d152,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D152, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d153,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D153, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d154,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D154, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d155,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D155, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d156,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D156, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d157,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D157, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d158,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D158, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d159,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D159, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d160,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D160, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d161,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D161, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d162,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D162, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d163,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D163, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d164,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D164, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d165,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D165, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d166,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D166, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d167,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D167, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d168,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D168, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d169,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D169, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d170,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D170, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d171,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D171, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d172,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D172, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d173,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D173, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d174,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D174, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d175,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D175, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d176,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D176, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d177,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D177, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d178,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D178, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d179,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D179, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d180,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D180, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d181,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D181, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d182,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D182, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d183,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D183, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d184,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D184, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d185,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D185, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d186,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D186, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d187,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D187, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d188,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D188, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d189,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D189, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d190,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D190, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d191,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D191, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d192,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D192, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d193,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D193, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d194,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D194, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d195,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D195, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d196,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D196, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d197,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D197, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d198,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D198, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d199,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D199, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d200,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D200, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d201,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D201, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d202,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D202, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d203,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D203, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d204,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D204, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d205,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D205, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d206,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D206, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d207,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D207, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d208,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D208, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d209,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D209, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d210,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D210, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d211,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D211, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d212,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D212, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d213,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D213, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d214,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D214, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d215,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D215, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d216,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D216, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d217,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D217, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d218,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D218, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d219,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D219, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d220,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D220, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d221,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D221, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d222,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D222, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d223,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D223, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d224,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D224, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d225,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D225, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d226,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D226, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d227,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D227, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d228,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D228, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d229,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D229, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d230,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D230, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d231,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D231, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d232,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D232, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d233,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D233, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d234,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D234, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d235,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D235, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d236,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D236, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d237,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D237, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d238,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D238, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d239,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D239, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d240,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D240, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d241,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D241, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d242,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D242, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d243,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D243, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d244,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D244, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d245,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D245, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d246,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D246, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d247,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D247, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d248,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D248, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d249,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D249, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d250,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D250, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d251,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D251, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d252,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D252, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d253,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D253, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d254,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D254, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d255,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D255, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d256,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D256, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d257,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D257, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d258,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D258, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d259,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D259, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d260,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D260, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d261,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D261, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d262,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D262, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d263,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D263, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d264,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D264, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d265,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D265, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d266,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D266, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d267,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D267, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d268,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D268, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d269,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D269, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d270,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D270, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d271,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D271, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d272,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D272, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d273,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D273, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d274,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D274, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d275,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D275, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d276,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D276, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d277,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D277, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d278,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D278, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d279,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D279, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d280,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D280, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d281,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D281, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d282,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D282, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d283,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D283, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d284,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D284, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d285,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D285, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d286,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D286, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d287,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D287, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d288,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D288, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d289,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D289, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d290,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D290, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d291,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D291, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d292,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D292, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d293,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D293, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d294,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D294, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d295,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D295, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d296,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D296, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d297,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D297, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d298,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D298, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d299,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D299, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d300,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D300, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d301,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D301, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d302,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D302, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d303,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D303, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d304,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D304, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d305,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D305, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d306,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D306, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d307,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D307, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d308,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D308, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d309,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D309, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d310,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D310, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d311,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D311, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d312,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D312, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d313,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D313, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d314,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D314, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d315,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D315, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d316,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D316, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d317,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D317, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d318,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D318, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d319,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D319, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d320,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D320, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d321,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D321, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d322,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D322, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d323,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D323, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d324,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D324, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d325,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D325, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d326,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D326, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d327,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D327, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d328,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D328, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d329,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D329, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d330,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D330, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d331,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D331, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d332,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D332, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d333,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D333, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d334,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D334, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d335,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D335, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d336,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D336, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d337,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D337, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d338,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D338, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d339,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D339, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d340,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D340, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d341,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D341, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d342,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D342, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d343,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D343, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d344,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D344, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d345,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D345, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d346,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D346, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d347,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D347, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d348,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D348, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d349,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D349, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d350,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D350, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d351,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D351, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d352,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D352, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d353,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D353, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d354,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D354, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d355,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D355, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d356,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D356, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d357,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D357, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d358,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D358, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d359,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D359, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d360,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D360, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d361,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D361, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d362,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D362, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d363,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D363, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d364,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D364, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d365,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D365, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d366,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D366, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d367,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D367, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d368,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D368, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d369,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D369, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d370,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D370, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d371,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D371, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d372,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D372, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d373,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D373, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d374,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D374, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d375,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D375, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d376,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D376, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d377,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D377, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d378,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D378, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d379,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D379, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d380,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D380, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d381,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D381, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d382,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D382, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d383,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D383, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d384,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D384, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d385,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D385, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d386,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D386, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d387,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D387, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d388,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D388, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d389,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D389, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d390,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D390, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d391,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D391, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d392,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D392, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d393,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D393, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d394,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D394, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d395,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D395, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d396,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D396, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d397,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D397, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d398,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D398, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d399,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D399, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d400,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D400, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d401,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D401, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d402,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D402, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d403,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D403, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d404,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D404, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d405,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D405, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d406,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D406, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d407,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D407, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d408,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D408, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d409,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D409, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d410,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D410, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d411,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D411, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d412,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D412, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d413,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D413, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d414,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D414, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d415,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D415, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d416,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D416, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d417,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D417, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d418,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D418, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d419,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D419, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d420,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D420, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d421,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D421, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d422,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D422, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d423,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D423, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d424,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D424, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d425,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D425, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d426,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D426, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d427,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D427, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d428,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D428, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d429,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D429, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d430,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D430, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d431,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D431, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d432,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D432, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d433,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D433, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d434,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D434, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d435,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D435, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d436,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D436, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d437,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D437, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d438,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D438, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d439,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D439, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d440,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D440, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d441,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D441, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d442,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D442, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d443,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D443, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d444,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D444, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d445,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D445, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d446,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D446, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d447,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D447, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d448,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D448, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d449,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D449, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d450,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D450, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d451,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D451, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d452,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D452, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d453,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D453, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d454,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D454, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d455,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D455, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d456,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D456, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d457,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D457, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d458,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D458, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d459,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D459, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d460,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D460, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d461,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D461, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d462,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D462, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d463,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D463, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d464,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D464, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d465,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D465, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d466,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D466, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d467,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D467, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d468,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D468, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d469,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D469, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d470,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D470, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d471,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D471, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d472,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D472, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d473,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D473, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d474,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D474, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d475,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D475, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d476,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D476, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d477,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D477, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d478,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D478, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d479,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D479, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d480,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D480, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d481,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D481, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d482,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D482, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d483,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D483, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d484,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D484, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d485,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D485, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d486,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D486, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d487,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D487, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d488,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D488, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d489,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D489, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d490,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D490, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d491,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D491, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d492,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D492, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d493,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D493, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d494,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D494, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d495,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D495, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d496,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D496, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d497,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D497, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d498,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D498, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d499,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D499, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d500,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D500, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d501,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D501, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d502,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D502, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d503,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D503, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d504,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D504, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d505,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D505, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d506,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D506, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d507,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D507, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d508,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D508, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d509,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D509, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d510,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D510, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d511,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D511, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d512,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D512, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d513,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D513, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d514,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D514, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d515,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D515, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d516,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D516, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d517,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D517, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d518,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D518, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d519,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D519, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d520,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D520, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d521,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D521, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d522,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D522, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d523,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D523, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d524,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D524, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d525,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D525, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d526,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D526, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d527,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D527, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d528,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D528, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d529,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D529, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d530,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D530, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d531,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D531, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d532,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D532, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d533,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D533, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d534,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D534, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d535,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D535, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d536,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D536, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d537,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D537, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d538,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D538, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d539,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D539, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d540,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D540, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d541,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D541, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d542,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D542, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d543,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D543, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d544,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D544, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d545,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D545, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d546,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D546, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d547,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D547, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d548,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D548, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d549,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D549, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d550,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D550, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d551,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D551, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d552,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D552, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d553,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D553, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d554,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D554, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d555,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D555, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d556,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D556, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d557,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D557, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d558,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D558, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d559,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D559, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d560,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D560, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d561,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D561, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d562,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D562, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d563,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D563, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d564,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D564, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d565,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D565, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d566,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D566, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d567,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D567, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d568,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D568, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d569,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D569, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d570,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D570, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d571,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D571, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d572,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D572, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d573,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D573, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d574,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D574, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d575,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D575, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d576,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D576, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d577,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D577, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d578,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D578, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d579,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D579, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d580,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D580, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d581,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D581, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d582,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D582, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d583,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D583, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d584,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D584, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d585,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D585, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d586,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D586, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d587,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D587, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d588,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D588, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d589,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D589, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d590,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D590, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d591,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D591, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d592,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D592, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d593,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D593, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d594,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D594, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d595,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D595, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d596,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D596, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d597,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D597, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d598,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D598, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d599,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D599, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d600,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D600, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d601,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D601, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d602,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D602, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d603,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D603, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d604,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D604, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d605,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D605, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d606,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D606, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d607,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D607, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d608,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D608, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d609,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D609, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d610,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D610, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d611,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D611, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d612,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D612, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d613,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D613, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d614,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D614, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d615,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D615, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d616,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D616, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d617,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D617, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d618,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D618, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d619,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D619, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d620,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D620, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d621,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D621, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d622,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D622, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d623,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D623, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d624,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D624, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d625,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D625, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d626,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D626, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d627,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D627, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d628,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D628, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d629,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D629, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d630,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D630, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d631,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D631, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d632,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D632, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d633,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D633, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d634,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D634, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d635,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D635, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d636,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D636, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d637,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D637, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d638,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D638, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d639,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D639, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d640,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D640, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d641,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D641, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d642,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D642, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d643,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D643, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d644,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D644, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d645,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D645, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d646,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D646, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d647,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D647, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d648,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D648, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d649,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D649, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d650,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D650, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d651,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D651, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d652,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D652, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d653,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D653, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d654,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D654, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d655,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D655, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d656,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D656, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d657,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D657, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d658,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D658, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d659,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D659, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d660,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D660, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d661,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D661, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d662,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D662, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d663,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D663, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d664,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D664, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d665,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D665, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d666,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D666, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d667,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D667, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d668,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D668, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d669,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D669, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d670,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D670, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d671,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D671, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d672,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D672, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d673,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D673, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d674,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D674, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d675,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D675, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d676,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D676, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d677,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D677, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d678,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D678, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d679,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D679, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d680,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D680, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d681,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D681, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d682,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D682, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d683,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D683, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d684,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D684, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d685,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D685, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d686,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D686, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d687,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D687, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d688,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D688, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d689,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D689, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d690,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D690, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d691,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D691, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d692,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D692, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d693,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D693, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d694,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D694, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d695,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D695, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d696,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D696, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d697,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D697, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d698,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D698, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d699,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D699, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d700,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D700, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d701,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D701, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d702,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D702, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d703,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D703, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d704,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D704, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d705,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D705, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d706,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D706, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d707,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D707, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d708,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D708, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d709,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D709, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d710,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D710, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d711,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D711, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d712,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D712, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d713,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D713, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d714,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D714, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d715,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D715, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d716,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D716, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d717,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D717, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d718,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D718, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d719,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D719, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d720,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D720, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d721,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D721, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d722,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D722, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d723,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D723, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d724,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D724, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d725,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D725, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d726,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D726, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d727,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D727, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d728,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D728, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d729,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D729, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d730,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D730, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d731,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D731, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d732,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D732, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d733,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D733, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d734,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D734, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d735,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D735, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d736,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D736, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d737,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D737, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d738,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D738, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d739,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D739, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d740,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D740, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d741,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D741, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d742,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D742, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d743,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D743, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d744,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D744, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d745,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D745, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d746,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D746, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d747,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D747, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d748,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D748, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d749,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D749, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d750,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D750, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d751,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D751, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d752,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D752, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d753,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D753, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d754,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D754, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d755,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D755, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d756,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D756, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d757,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D757, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d758,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D758, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d759,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D759, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d760,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D760, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d761,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D761, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d762,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D762, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d763,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D763, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d764,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D764, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d765,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D765, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d766,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D766, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d767,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D767, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d768,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D768, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d769,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D769, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d770,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D770, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d771,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D771, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d772,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D772, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d773,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D773, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d774,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D774, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d775,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D775, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d776,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D776, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d777,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D777, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d778,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D778, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d779,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D779, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d780,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D780, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d781,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D781, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d782,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D782, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d783,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D783, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d784,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D784, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d785,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D785, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d786,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D786, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d787,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D787, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d788,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D788, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d789,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D789, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d790,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D790, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d791,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D791, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d792,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D792, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d793,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D793, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d794,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D794, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d795,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D795, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d796,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D796, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d797,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D797, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d798,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D798, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d799,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D799, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d800,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D800, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d801,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D801, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d802,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D802, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d803,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D803, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d804,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D804, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d805,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D805, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d806,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D806, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d807,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D807, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d808,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D808, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d809,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D809, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d810,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D810, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d811,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D811, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d812,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D812, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d813,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D813, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d814,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D814, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d815,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D815, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d816,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D816, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d817,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D817, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d818,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D818, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d819,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D819, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d820,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D820, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d821,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D821, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d822,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D822, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d823,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D823, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d824,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D824, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d825,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D825, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d826,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D826, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d827,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D827, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d828,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D828, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d829,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D829, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d830,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D830, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d831,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D831, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d832,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D832, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d833,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D833, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d834,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D834, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d835,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D835, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d836,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D836, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d837,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D837, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d838,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D838, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d839,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D839, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d840,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D840, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d841,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D841, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d842,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D842, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d843,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D843, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d844,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D844, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d845,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D845, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d846,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D846, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d847,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D847, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d848,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D848, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d849,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D849, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d850,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D850, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d851,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D851, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d852,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D852, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d853,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D853, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d854,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D854, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d855,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D855, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d856,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D856, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d857,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D857, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d858,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D858, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d859,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D859, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d860,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D860, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d861,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D861, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d862,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D862, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d863,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D863, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d864,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D864, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d865,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D865, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d866,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D866, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d867,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D867, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d868,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D868, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d869,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D869, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d870,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D870, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d871,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D871, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d872,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D872, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d873,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D873, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d874,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D874, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d875,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D875, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d876,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D876, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d877,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D877, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d878,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D878, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d879,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D879, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d880,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D880, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d881,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D881, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d882,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D882, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d883,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D883, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d884,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D884, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d885,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D885, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d886,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D886, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d887,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D887, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d888,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D888, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d889,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D889, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d890,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D890, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d891,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D891, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d892,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D892, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d893,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D893, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d894,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D894, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d895,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D895, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d896,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D896, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d897,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D897, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d898,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D898, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d899,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D899, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d900,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D900, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d901,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D901, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d902,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D902, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d903,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D903, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d904,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D904, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d905,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D905, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d906,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D906, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d907,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D907, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d908,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D908, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d909,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D909, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d910,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D910, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d911,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D911, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d912,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D912, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d913,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D913, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d914,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D914, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d915,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D915, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d916,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D916, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d917,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D917, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d918,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D918, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d919,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D919, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d920,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D920, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d921,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D921, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d922,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D922, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d923,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D923, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d924,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D924, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d925,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D925, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d926,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D926, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d927,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D927, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d928,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D928, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d929,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D929, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d930,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D930, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d931,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D931, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d932,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D932, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d933,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D933, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d934,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D934, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d935,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D935, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d936,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D936, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d937,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D937, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d938,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D938, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d939,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D939, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d940,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D940, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d941,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D941, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d942,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D942, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d943,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D943, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d944,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D944, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d945,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D945, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d946,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D946, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d947,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D947, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d948,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D948, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d949,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D949, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d950,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D950, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d951,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D951, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d952,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D952, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d953,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D953, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d954,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D954, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d955,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D955, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d956,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D956, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d957,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D957, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d958,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D958, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d959,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D959, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d960,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D960, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d961,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D961, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d962,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D962, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d963,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D963, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d964,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D964, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d965,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D965, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d966,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D966, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d967,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D967, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d968,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D968, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d969,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D969, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d970,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D970, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d971,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D971, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d972,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D972, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d973,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D973, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d974,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D974, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d975,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D975, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d976,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D976, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d977,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D977, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d978,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D978, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d979,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D979, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d980,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D980, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d981,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D981, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d982,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D982, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d983,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D983, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d984,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D984, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d985,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D985, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d986,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D986, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d987,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D987, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d988,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D988, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d989,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D989, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d990,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D990, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d991,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D991, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d992,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D992, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d993,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D993, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d994,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D994, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d995,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D995, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d996,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D996, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d997,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D997, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d998,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D998, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d999,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D999, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1000,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1000, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1001,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1001, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1002,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1002, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1003,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1003, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1004,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1004, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1005,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1005, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1006,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1006, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1007,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1007, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1008,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1008, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1009,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1009, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1010,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1010, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1011,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1011, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1012,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1012, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1013,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1013, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1014,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1014, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1015,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1015, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1016,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1016, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1017,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1017, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1018,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1018, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1019,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1019, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1020,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1020, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1021,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1021, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1022,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1022, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1023,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1023, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1024,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1024, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1025,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1025, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1026,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1026, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1027,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1027, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1028,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1028, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1029,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1029, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1030,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1030, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1031,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1031, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1032,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1032, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1033,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1033, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1034,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1034, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1035,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1035, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1036,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1036, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1037,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1037, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1038,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1038, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1039,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1039, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1040,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1040, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1041,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1041, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1042,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1042, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1043,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1043, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1044,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1044, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1045,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1045, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1046,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1046, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1047,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1047, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1048,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1048, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1049,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1049, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1050,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1050, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1051,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1051, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1052,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1052, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1053,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1053, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1054,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1054, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1055,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1055, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1056,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1056, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1057,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1057, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1058,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1058, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1059,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1059, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1060,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1060, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1061,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1061, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1062,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1062, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1063,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1063, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1064,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1064, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1065,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1065, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1066,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1066, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1067,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1067, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1068,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1068, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1069,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1069, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1070,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1070, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1071,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1071, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1072,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1072, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1073,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1073, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1074,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1074, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1075,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1075, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1076,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1076, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1077,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1077, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1078,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1078, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1079,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1079, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1080,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1080, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1081,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1081, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1082,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1082, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1083,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1083, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1084,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1084, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1085,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1085, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1086,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1086, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1087,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1087, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1088,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1088, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1089,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1089, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1090,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1090, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1091,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1091, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1092,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1092, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1093,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1093, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1094,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1094, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1095,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1095, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1096,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1096, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1097,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1097, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1098,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1098, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1099,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1099, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1100,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1100, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1101,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1101, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1102,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1102, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1103,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1103, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1104,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1104, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1105,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1105, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1106,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1106, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1107,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1107, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1108,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1108, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1109,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1109, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1110,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1110, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1111,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1111, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1112,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1112, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1113,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1113, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1114,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1114, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1115,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1115, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1116,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1116, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1117,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1117, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1118,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1118, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1119,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1119, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1120,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1120, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1121,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1121, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1122,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1122, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1123,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1123, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1124,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1124, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1125,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1125, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1126,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1126, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1127,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1127, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1128,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1128, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1129,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1129, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1130,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1130, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1131,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1131, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1132,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1132, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1133,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1133, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1134,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1134, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1135,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1135, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1136,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1136, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1137,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1137, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1138,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1138, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1139,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1139, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1140,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1140, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1141,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1141, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1142,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1142, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1143,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1143, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1144,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1144, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1145,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1145, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1146,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1146, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1147,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1147, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1148,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1148, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1149,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1149, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1150,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1150, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1151,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1151, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1152,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1152, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1153,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1153, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1154,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1154, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1155,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1155, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1156,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1156, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1157,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1157, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1158,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1158, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1159,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1159, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1160,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1160, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1161,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1161, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1162,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1162, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1163,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1163, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1164,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1164, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1165,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1165, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1166,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1166, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1167,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1167, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1168,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1168, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1169,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1169, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1170,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1170, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1171,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1171, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1172,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1172, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1173,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1173, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1174,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1174, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1175,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1175, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1176,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1176, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1177,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1177, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1178,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1178, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1179,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1179, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1180,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1180, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1181,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1181, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1182,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1182, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1183,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1183, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1184,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1184, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1185,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1185, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1186,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1186, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1187,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1187, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1188,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1188, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1189,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1189, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1190,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1190, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1191,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1191, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1192,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1192, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1193,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1193, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1194,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1194, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1195,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1195, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1196,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1196, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1197,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1197, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1198,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1198, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1199,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1199, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1200,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1200, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1201,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1201, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1202,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1202, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1203,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1203, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1204,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1204, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1205,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1205, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1206,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1206, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1207,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1207, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1208,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1208, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1209,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1209, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1210,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1210, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1211,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1211, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1212,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1212, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1213,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1213, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1214,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1214, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1215,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1215, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1216,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1216, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1217,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1217, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1218,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1218, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1219,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1219, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1220,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1220, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1221,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1221, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1222,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1222, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1223,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1223, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1224,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1224, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1225,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1225, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1226,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1226, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1227,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1227, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1228,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1228, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1229,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1229, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1230,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1230, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1231,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1231, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1232,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1232, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1233,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1233, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1234,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1234, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1235,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1235, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1236,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1236, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1237,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1237, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1238,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1238, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1239,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1239, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1240,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1240, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1241,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1241, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1242,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1242, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1243,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1243, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1244,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1244, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1245,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1245, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1246,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1246, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1247,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1247, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1248,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1248, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1249,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1249, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1250,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1250, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1251,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1251, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1252,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1252, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1253,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1253, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1254,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1254, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1255,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1255, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1256,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1256, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1257,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1257, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1258,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1258, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1259,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1259, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1260,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1260, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1261,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1261, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1262,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1262, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1263,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1263, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1264,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1264, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1265,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1265, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1266,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1266, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1267,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1267, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1268,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1268, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1269,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1269, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1270,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1270, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1271,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1271, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1272,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1272, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1273,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1273, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1274,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1274, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1275,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1275, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1276,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1276, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1277,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1277, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1278,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1278, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1279,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1279, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1280,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1280, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1281,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1281, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1282,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1282, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1283,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1283, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1284,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1284, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1285,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1285, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1286,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1286, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1287,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1287, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1288,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1288, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1289,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1289, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1290,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1290, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1291,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1291, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1292,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1292, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1293,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1293, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1294,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1294, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1295,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1295, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1296,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1296, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1297,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1297, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1298,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1298, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1299,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1299, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1300,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1300, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1301,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1301, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1302,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1302, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1303,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1303, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1304,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1304, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1305,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1305, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1306,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1306, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1307,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1307, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1308,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1308, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1309,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1309, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1310,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1310, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1311,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1311, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1312,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1312, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1313,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1313, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1314,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1314, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1315,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1315, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1316,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1316, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1317,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1317, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1318,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1318, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1319,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1319, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1320,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1320, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1321,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1321, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1322,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1322, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1323,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1323, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1324,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1324, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1325,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1325, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1326,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1326, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1327,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1327, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1328,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1328, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1329,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1329, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1330,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1330, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1331,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1331, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1332,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1332, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1333,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1333, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1334,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1334, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1335,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1335, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1336,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1336, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1337,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1337, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1338,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1338, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1339,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1339, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1340,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1340, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1341,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1341, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1342,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1342, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1343,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1343, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1344,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1344, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1345,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1345, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1346,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1346, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1347,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1347, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1348,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1348, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1349,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1349, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1350,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1350, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1351,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1351, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1352,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1352, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1353,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1353, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1354,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1354, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1355,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1355, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1356,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1356, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1357,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1357, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1358,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1358, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1359,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1359, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1360,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1360, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1361,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1361, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1362,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1362, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1363,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1363, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1364,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1364, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1365,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1365, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1366,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1366, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1367,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1367, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1368,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1368, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1369,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1369, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1370,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1370, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1371,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1371, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1372,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1372, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1373,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1373, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1374,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1374, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1375,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1375, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1376,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1376, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1377,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1377, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1378,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1378, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1379,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1379, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1380,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1380, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1381,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1381, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1382,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1382, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1383,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1383, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1384,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1384, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1385,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1385, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1386,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1386, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1387,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1387, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1388,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1388, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1389,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1389, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1390,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1390, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1391,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1391, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1392,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1392, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1393,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1393, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1394,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1394, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1395,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1395, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1396,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1396, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1397,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1397, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1398,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1398, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1399,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1399, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1400,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1400, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1401,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1401, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1402,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1402, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1403,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1403, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1404,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1404, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1405,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1405, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1406,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1406, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1407,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1407, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1408,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1408, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1409,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1409, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1410,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1410, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1411,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1411, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1412,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1412, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1413,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1413, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1414,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1414, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1415,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1415, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1416,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1416, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1417,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1417, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1418,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1418, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1419,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1419, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1420,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1420, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1421,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1421, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1422,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1422, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1423,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1423, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1424,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1424, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1425,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1425, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1426,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1426, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1427,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1427, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1428,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1428, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1429,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1429, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1430,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1430, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1431,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1431, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1432,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1432, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1433,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1433, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1434,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1434, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1435,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1435, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1436,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1436, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1437,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1437, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1438,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1438, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1439,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1439, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1440,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1440, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1441,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1441, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1442,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1442, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1443,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1443, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1444,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1444, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1445,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1445, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1446,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1446, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1447,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1447, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1448,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1448, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1449,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1449, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1450,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1450, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1451,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1451, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1452,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1452, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1453,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1453, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1454,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1454, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1455,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1455, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1456,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1456, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1457,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1457, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1458,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1458, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1459,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1459, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1460,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1460, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1461,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1461, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1462,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1462, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1463,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1463, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1464,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1464, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1465,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1465, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1466,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1466, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1467,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1467, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1468,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1468, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1469,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1469, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1470,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1470, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1471,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1471, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1472,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1472, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1473,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1473, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1474,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1474, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1475,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1475, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1476,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1476, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1477,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1477, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1478,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1478, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1479,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1479, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1480,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1480, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1481,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1481, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1482,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1482, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1483,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1483, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1484,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1484, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1485,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1485, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1486,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1486, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1487,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1487, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1488,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1488, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1489,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1489, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1490,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1490, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1491,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1491, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1492,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1492, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1493,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1493, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1494,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1494, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1495,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1495, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1496,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1496, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1497,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1497, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1498,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1498, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1499,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1499, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1500,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1500, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1501,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1501, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1502,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1502, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1503,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1503, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1504,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1504, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1505,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1505, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1506,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1506, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1507,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1507, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1508,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1508, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1509,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1509, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1510,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1510, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1511,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1511, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1512,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1512, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1513,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1513, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1514,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1514, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1515,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1515, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1516,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1516, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1517,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1517, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1518,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1518, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1519,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1519, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1520,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1520, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1521,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1521, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1522,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1522, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1523,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1523, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1524,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1524, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1525,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1525, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1526,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1526, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1527,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1527, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1528,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1528, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1529,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1529, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1530,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1530, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1531,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1531, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1532,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1532, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1533,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1533, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1534,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1534, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1535,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1535, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1536,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1536, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1537,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1537, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1538,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1538, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1539,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1539, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1540,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1540, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1541,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1541, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1542,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1542, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1543,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1543, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1544,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1544, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1545,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1545, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1546,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1546, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1547,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1547, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1548,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1548, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1549,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1549, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1550,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1550, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1551,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1551, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1552,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1552, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1553,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1553, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1554,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1554, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1555,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1555, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1556,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1556, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1557,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1557, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1558,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1558, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1559,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1559, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1560,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1560, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1561,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1561, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1562,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1562, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1563,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1563, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1564,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1564, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1565,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1565, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1566,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1566, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1567,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1567, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1568,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1568, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1569,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1569, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1570,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1570, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1571,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1571, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1572,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1572, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1573,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1573, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1574,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1574, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1575,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1575, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1576,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1576, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1577,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1577, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1578,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1578, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1579,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1579, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1580,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1580, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1581,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1581, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1582,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1582, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1583,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1583, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1584,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1584, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1585,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1585, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1586,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1586, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1587,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1587, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1588,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1588, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1589,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1589, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1590,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1590, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1591,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1591, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1592,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1592, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1593,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1593, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1594,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1594, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1595,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1595, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1596,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1596, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1597,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1597, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1598,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1598, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1599,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1599, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1600,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1600, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1601,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1601, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1602,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1602, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1603,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1603, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1604,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1604, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1605,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1605, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1606,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1606, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1607,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1607, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1608,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1608, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1609,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1609, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1610,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1610, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1611,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1611, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1612,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1612, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1613,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1613, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1614,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1614, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1615,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1615, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1616,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1616, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1617,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1617, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1618,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1618, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1619,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1619, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1620,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1620, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1621,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1621, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1622,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1622, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1623,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1623, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1624,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1624, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1625,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1625, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1626,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1626, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1627,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1627, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1628,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1628, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1629,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1629, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1630,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1630, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1631,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1631, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1632,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1632, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1633,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1633, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1634,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1634, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1635,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1635, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1636,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1636, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1637,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1637, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1638,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1638, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1639,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1639, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1640,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1640, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1641,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1641, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1642,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1642, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1643,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1643, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1644,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1644, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1645,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1645, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1646,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1646, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1647,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1647, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1648,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1648, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1649,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1649, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1650,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1650, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1651,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1651, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1652,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1652, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1653,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1653, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1654,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1654, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1655,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1655, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1656,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1656, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1657,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1657, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1658,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1658, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1659,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1659, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1660,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1660, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1661,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1661, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1662,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1662, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1663,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1663, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1664,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1664, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1665,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1665, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1666,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1666, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1667,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1667, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1668,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1668, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1669,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1669, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1670,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1670, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1671,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1671, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1672,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1672, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1673,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1673, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1674,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1674, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1675,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1675, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1676,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1676, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1677,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1677, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1678,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1678, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1679,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1679, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1680,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1680, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1681,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1681, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1682,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1682, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1683,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1683, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1684,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1684, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1685,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1685, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1686,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1686, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1687,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1687, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1688,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1688, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1689,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1689, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1690,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1690, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1691,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1691, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1692,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1692, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1693,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1693, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1694,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1694, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1695,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1695, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1696,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1696, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1697,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1697, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1698,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1698, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1699,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1699, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1700,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1700, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1701,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1701, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1702,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1702, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1703,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1703, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1704,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1704, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1705,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1705, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1706,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1706, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1707,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1707, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1708,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1708, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1709,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1709, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1710,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1710, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1711,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1711, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1712,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1712, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1713,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1713, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1714,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1714, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1715,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1715, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1716,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1716, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1717,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1717, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1718,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1718, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1719,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1719, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1720,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1720, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1721,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1721, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1722,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1722, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1723,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1723, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1724,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1724, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1725,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1725, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1726,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1726, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1727,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1727, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1728,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1728, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1729,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1729, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1730,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1730, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1731,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1731, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1732,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1732, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1733,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1733, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1734,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1734, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1735,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1735, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1736,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1736, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1737,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1737, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1738,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1738, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1739,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1739, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1740,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1740, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1741,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1741, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1742,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1742, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1743,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1743, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1744,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1744, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1745,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1745, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1746,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1746, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1747,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1747, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1748,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1748, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1749,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1749, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1750,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1750, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1751,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1751, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1752,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1752, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1753,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1753, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1754,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1754, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1755,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1755, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1756,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1756, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1757,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1757, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1758,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1758, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1759,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1759, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1760,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1760, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1761,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1761, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1762,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1762, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1763,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1763, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1764,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1764, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1765,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1765, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1766,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1766, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1767,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1767, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1768,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1768, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1769,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1769, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1770,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1770, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1771,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1771, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1772,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1772, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1773,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1773, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1774,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1774, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1775,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1775, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1776,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1776, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1777,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1777, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1778,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1778, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1779,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1779, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1780,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1780, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1781,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1781, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1782,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1782, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1783,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1783, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1784,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1784, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1785,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1785, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1786,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1786, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1787,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1787, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1788,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1788, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1789,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1789, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1790,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1790, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1791,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1791, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1792,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1792, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1793,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1793, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1794,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1794, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1795,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1795, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1796,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1796, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1797,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1797, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1798,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1798, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1799,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1799, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1800,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1800, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1801,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1801, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1802,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1802, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1803,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1803, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1804,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1804, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1805,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1805, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1806,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1806, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1807,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1807, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1808,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1808, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1809,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1809, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1810,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1810, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1811,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1811, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1812,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1812, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1813,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1813, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1814,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1814, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1815,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1815, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1816,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1816, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1817,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1817, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1818,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1818, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1819,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1819, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1820,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1820, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1821,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1821, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1822,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1822, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1823,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1823, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1824,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1824, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1825,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1825, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1826,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1826, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1827,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1827, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1828,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1828, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1829,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1829, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1830,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1830, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1831,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1831, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1832,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1832, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1833,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1833, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1834,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1834, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1835,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1835, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1836,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1836, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1837,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1837, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1838,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1838, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1839,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1839, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1840,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1840, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1841,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1841, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1842,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1842, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1843,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1843, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1844,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1844, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1845,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1845, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1846,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1846, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1847,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1847, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1848,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1848, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1849,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1849, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1850,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1850, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1851,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1851, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1852,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1852, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1853,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1853, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1854,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1854, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1855,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1855, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1856,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1856, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1857,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1857, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1858,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1858, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1859,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1859, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1860,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1860, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1861,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1861, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1862,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1862, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1863,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1863, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1864,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1864, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1865,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1865, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1866,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1866, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1867,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1867, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1868,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1868, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1869,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1869, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1870,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1870, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1871,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1871, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1872,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1872, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1873,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1873, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1874,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1874, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1875,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1875, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1876,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1876, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1877,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1877, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1878,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1878, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1879,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1879, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1880,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1880, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1881,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1881, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1882,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1882, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1883,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1883, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1884,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1884, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1885,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1885, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1886,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1886, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1887,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1887, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1888,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1888, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1889,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1889, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1890,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1890, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1891,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1891, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1892,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1892, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1893,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1893, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1894,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1894, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1895,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1895, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1896,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1896, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1897,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1897, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1898,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1898, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1899,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1899, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1900,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1900, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1901,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1901, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1902,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1902, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1903,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1903, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1904,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1904, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1905,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1905, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1906,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1906, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1907,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1907, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1908,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1908, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1909,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1909, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1910,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1910, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1911,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1911, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1912,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1912, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1913,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1913, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1914,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1914, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1915,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1915, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1916,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1916, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1917,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1917, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1918,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1918, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1919,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1919, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1920,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1920, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1921,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1921, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1922,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1922, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1923,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1923, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1924,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1924, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1925,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1925, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1926,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1926, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1927,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1927, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1928,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1928, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1929,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1929, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1930,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1930, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1931,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1931, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1932,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1932, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1933,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1933, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1934,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1934, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1935,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1935, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1936,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1936, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1937,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1937, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1938,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1938, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1939,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1939, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1940,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1940, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1941,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1941, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1942,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1942, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1943,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1943, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1944,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1944, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1945,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1945, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1946,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1946, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1947,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1947, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1948,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1948, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1949,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1949, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1950,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1950, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1951,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1951, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1952,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1952, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1953,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1953, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1954,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1954, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1955,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1955, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1956,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1956, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1957,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1957, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1958,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1958, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1959,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1959, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1960,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1960, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1961,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1961, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1962,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1962, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1963,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1963, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1964,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1964, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1965,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1965, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1966,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1966, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1967,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1967, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1968,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1968, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1969,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1969, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1970,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1970, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1971,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1971, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1972,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1972, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1973,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1973, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1974,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1974, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1975,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1975, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1976,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1976, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1977,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1977, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1978,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1978, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1979,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1979, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1980,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1980, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1981,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1981, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1982,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1982, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1983,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1983, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1984,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1984, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1985,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1985, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1986,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1986, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1987,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1987, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1988,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1988, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1989,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1989, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1990,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1990, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1991,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1991, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1992,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1992, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1993,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1993, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1994,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1994, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1995,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1995, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1996,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1996, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1997,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1997, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1998,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1998, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d1999,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1999, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d2000,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2000, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d2001,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2001, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d2002,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2002, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d2003,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2003, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d2004,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2004, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d2005,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2005, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d2006,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2006, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d2007,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2007, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d2008,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2008, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d2009,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2009, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d2010,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2010, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d2011,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2011, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d2012,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2012, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d2013,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2013, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d2014,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2014, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d2015,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2015, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d2016,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2016, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d2017,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2017, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d2018,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2018, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d2019,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2019, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d2020,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2020, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d2021,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2021, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d2022,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2022, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d2023,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2023, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d2024,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2024, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d2025,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2025, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d2026,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2026, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d2027,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2027, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d2028,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2028, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d2029,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2029, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d2030,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2030, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d2031,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2031, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d2032,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2032, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d2033,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2033, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d2034,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2034, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d2035,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2035, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d2036,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2036, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d2037,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2037, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d2038,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2038, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d2039,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2039, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d2040,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2040, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d2041,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2041, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d2042,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2042, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d2043,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2043, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d2044,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2044, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d2045,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2045, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d2046,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2046, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     

       begin//{ 
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================
         `payload_generate('h0,'d2047,'h1,local_fmt_type);
         
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2047, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         fmt_type    == local_fmt_type    ;
                                                                         direction   == 1'b1              ;             
                                                                                              })
                    
         end//}     


  
join_none
wait fork;	
