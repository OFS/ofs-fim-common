// Copyright 2022 Intel Corporation
// SPDX-License-Identifier: MIT
//
// Create Date  : Feb 2021
// Module Name  : protocol_checker_csr.sv
// Project      : OFS
// -----------------------------------------------------------------------------
//
// ***************************************************************************


// BEGIN TEMPLATE
//
// *******************************************************
// *** WARNING!! ** WARNING!! ** WARNING!! ** WARNING!!***
// ***             DO NOT EDIT THIS FILE!!             ***
// *******************************************************
// This file is automatically generated from the files:
// ./protocol_checker_csrs.ini and ./protocol_checker_csr_template.sv using the perl
// program mk_reg_def.pl. Modify one of these files if you wish to make a change to
// this file.
//
// The mk_cfg_module_64.pl script generates these files:
//         Register Block RTL (this file) ./protocol_checker_csr.sv
//         The Register Specification     ./protocol_checker_csr_spec.html
//
// The input files used are:
//         register definition file       ./protocol_checker_csrs.ini
//         Register Block Template        ./protocol_checker_csr_template.sv
//         The perl script                ../../../tools/mk_csr_module\mk_cfg_module_64.pl
//
module  protocol_checker_csr
  import ofs_csr_pkg::*;
   import prtcl_chkr_pkg::*;
   #(parameter HI_ADDR_BIT = 11     )(
       input        clk_csr,
       input        rst_n_csr,
       input        pwr_good_csr_clk_n,
       input        pwr_good_clk_n,
       input        clk,
       input        rst_n,
       input        i_blocking_traffic,
       ofs_fim_axi_lite_if.slave csr_lite_if,
       t_prtcl_chkr_err_vector i_error_vector,
       t_mmio_timeout_hdr_info i_mmio_timeout_info,
       output logic o_clear_errors
       
       
       // BELOW IS A KEY PHRASE THE mk_cfg_module_64.pl
       // KEYS ON. DO NOT DELETE.
       // ***************************************
       // Start Auto generated input port list (string key for mk_cfg_module_64.pl)
       // ***************************************
   ,input logic[10:00] i_vf_num_load_data                  // load data for register  0x010 afu_intf_error            bits 28:18 (vf_num)
   ,input logic        i_tx_hdr_is_pu_mode_load_data       // load data for register  0x030 mmio_immediate_frozen_reg bit  01    (tx_hdr_is_pu_mode)
   ,input logic        i_mmio_immediate_frozen_load_data   // load data for register  0x030 mmio_immediate_frozen_reg bit  00    (mmio_immediate_frozen)
   ,input logic[63:00] i_tx_header_error_255_192_load_data // load data for register  0x038 mmio_tx_header_error_255_192 bits 63:00 (tx_header_error_255_192)
   ,input logic[63:00] i_tx_header_error_191_128_load_data // load data for register  0x040 mmio_tx_header_error_191_128 bits 63:00 (tx_header_error_191_128)
   ,input logic[63:00] i_tx_header_error_127_64_load_data  // load data for register  0x048 mmio_tx_header_error_127_64 bits 63:00 (tx_header_error_127_64)
   ,input logic[63:00] i_tx_header_error_63_00_load_data   // load data for register  0x050 mmio_tx_header_error_63_00 bits 63:00 (tx_header_error_63_00)
       
       // BELOW IS A KEY PHRASE THE mk_cfg_module_64.pl
       // KEYS ON. DO NOT DELETE.
       // ***************************************
       // Start Auto generated output port list (string key for mk_cfg_module_64.pl)
       // ***************************************
       );
   
   // BELOW IS A KEY PHRASE THE mk_cfg_module_64.pl
   // KEYS ON. DO NOT DELETE.
   // ***************************************
   // Start Auto generated reg and wire decls (string key for mk_cfg_module_64.pl)
   // ***************************************
   logic   decode_11_8_00;
   logic   decode_11_8_01;
   logic   decode_11_8_02;
   logic   decode_11_8_03;
   logic   decode_11_8_04;
   logic   decode_11_8_05;
   logic   decode_11_8_06;
   logic   decode_11_8_07;
   logic   decode_11_8_08;
   logic   decode_11_8_09;
   logic   decode_11_8_10;
   logic   decode_11_8_11;
   logic   decode_11_8_12;
   logic   decode_11_8_13;
   logic   decode_11_8_14;
   logic   decode_11_8_15;

   // ******************************************************
   // Register 0x000 afu_intf_dfh
   // ******************************************************
   logic [63:00] afu_intf_dfh_wire;                       // Register 0x000
   logic [03:00] feature_type_reg;                        // bit(s) 63:60
   logic         eol_reg;                                 // bit(s) 40:40
   logic [23:00] next_dfh_byte_offset_reg;                // bit(s) 39:16
   logic [03:00] feature_rev_reg;                         // bit(s) 15:12
   logic [11:00] feature_id_reg;                          // bit(s) 11:00


   // ******************************************************
   // Register 0x008 afu_intf_scratchpad
   // ******************************************************
   logic [63:00] afu_intf_scratchpad_wire;                // Register 0x008
   logic [63:00] scratchpad_reg;                          // bit(s) 63:00


   // ******************************************************
   // Register 0x010 afu_intf_error
   // ******************************************************
   logic [63:00] afu_intf_error_wire;                     // Register 0x010
   logic         blocking_traffic_reg;                    // bit(s) 31:31
   logic [10:00] vf_num_reg;                              // bit(s) 28:18
   logic         vf_flr_access_reg;                       // bit(s) 17:17
   logic         malformed_tlp_err_reg;                   // bit(s) 14:14
   logic         max_payload_err_reg;                     // bit(s) 13:13
   logic         max_read_req_size_err_reg;               // bit(s) 12:12
   logic         max_tag_err_reg;                         // bit(s) 11:11
   logic         unexp_mmio_rsp_err_reg;                  // bit(s) 08:08
   logic         mmio_timeout_err_reg;                    // bit(s) 07:07
   logic         mmio_data_payload_overrun_err_reg;       // bit(s) 04:04
   logic         mmio_insufficient_data_err_reg;          // bit(s) 03:03
   logic         tx_mwr_data_payload_overrun_err_reg;     // bit(s) 02:02
   logic         tx_mwr_insufficient_data_err_reg;        // bit(s) 01:01


   // ******************************************************
   // Register 0x018 afu_intf_first_error
   // ******************************************************
   logic [63:00] afu_intf_first_error_wire;               // Register 0x018
   logic [10:00] vf_num_ferr_reg;                         // bit(s) 28:18
   logic         vf_flr_access_ferr_reg;                  // bit(s) 17:17
   logic         malformed_tlp_ferr_reg;                  // bit(s) 14:14
   logic         max_payload_ferr_reg;                    // bit(s) 13:13
   logic         max_read_req_size_ferr_reg;              // bit(s) 12:12
   logic         max_tag_ferr_reg;                        // bit(s) 11:11
   logic         unexp_mmio_rsp_ferr_reg;                 // bit(s) 08:08
   logic         mmio_timeout_ferr_reg;                   // bit(s) 07:07
   logic         mmio_data_payload_overrun_ferr_reg;      // bit(s) 04:04
   logic         mmio_insufficient_data_ferr_reg;         // bit(s) 03:03
   logic         tx_mwr_data_payload_overrun_ferr_reg;    // bit(s) 02:02
   logic         tx_mwr_insufficient_data_ferr_reg;       // bit(s) 01:01


   // ******************************************************
   // Register 0x020 mmio_timeout_addr
   // ******************************************************
   logic [63:00] mmio_timeout_addr_wire;                  // Register 0x020
   logic [31:00] mmio_timeout_addr_reg;                   // bit(s) 31:00


   // ******************************************************
   // Register 0x028 mmio_timeout_info
   // ******************************************************
   logic [63:00] mmio_timeout_info_wire;                  // Register 0x028
   logic         timeout_regs_frozen_reg;                 // bit(s) 63:63
   logic [07:00] mmio_timeout_tag_reg;                    // bit(s) 35:28
   logic [09:00] mmio_timeout_dw0_len_reg;                // bit(s) 25:16
   logic [15:00] mmio_timeout_requester_id_reg;           // bit(s) 15:00


   // ******************************************************
   // Register 0x030 mmio_immediate_frozen_reg
   // ******************************************************
   logic [63:00] mmio_immediate_frozen_reg_wire;          // Register 0x030
   logic         tx_hdr_is_pu_mode_reg;                   // bit(s) 01:01
   logic         mmio_immediate_frozen_reg;               // bit(s) 00:00


   // ******************************************************
   // Register 0x038 mmio_tx_header_error_255_192
   // ******************************************************
   logic [63:00] mmio_tx_header_error_255_192_wire;       // Register 0x038
   logic [63:00] tx_header_error_255_192_reg;             // bit(s) 63:00


   // ******************************************************
   // Register 0x040 mmio_tx_header_error_191_128
   // ******************************************************
   logic [63:00] mmio_tx_header_error_191_128_wire;       // Register 0x040
   logic [63:00] tx_header_error_191_128_reg;             // bit(s) 63:00


   // ******************************************************
   // Register 0x048 mmio_tx_header_error_127_64
   // ******************************************************
   logic [63:00] mmio_tx_header_error_127_64_wire;        // Register 0x048
   logic [63:00] tx_header_error_127_64_reg;              // bit(s) 63:00


   // ******************************************************
   // Register 0x050 mmio_tx_header_error_63_00
   // ******************************************************
   logic [63:00] mmio_tx_header_error_63_00_wire;         // Register 0x050
   logic [63:00] tx_header_error_63_00_reg;               // bit(s) 63:00

   logic         rd_or_wr_r2;

   // *****************************************************
   // Logic declairs for the 8 bit "register" decode nets.
   // *****************************************************
   logic         afu_intf_dfh_en_r3;
   logic         afu_intf_scratchpad_en_r3;
   logic         afu_intf_error_en_r3;
   logic         afu_intf_first_error_en_r3;
   logic         mmio_timeout_addr_en_r3;
   logic         mmio_timeout_info_en_r3;
   logic         mmio_immediate_frozen_reg_en_r3;
   logic         mmio_tx_header_error_255_192_en_r3;
   logic         mmio_tx_header_error_191_128_en_r3;
   logic         mmio_tx_header_error_127_64_en_r3;
   logic         mmio_tx_header_error_63_00_en_r3;
   logic [63:00] csr_decode_mux_r4;
   // ******************************************************
   // *declair logics that are terms but not ports.
   // ******************************************************
  logic          set_malformed_tlp_err; // set term for register 0x010 afu_intf_error bit(s) 14:14 (malformed_tlp_err)
  logic          set_max_payload_err; // set term for register 0x010 afu_intf_error bit(s) 13:13 (max_payload_err)
  logic          set_max_read_req_size_err; // set term for register 0x010 afu_intf_error bit(s) 12:12 (max_read_req_size_err)
  logic          set_max_tag_err; // set term for register 0x010 afu_intf_error bit(s) 11:11 (max_tag_err)
  logic          set_unexp_mmio_rsp_err; // set term for register 0x010 afu_intf_error bit(s) 08:08 (unexp_mmio_rsp_err)
  logic          set_mmio_timeout_err; // set term for register 0x010 afu_intf_error bit(s) 07:07 (mmio_timeout_err)
  logic          set_mmio_data_payload_overrun_err; // set term for register 0x010 afu_intf_error bit(s) 04:04 (mmio_data_payload_overrun_err)
  logic          set_mmio_insufficient_data_err; // set term for register 0x010 afu_intf_error bit(s) 03:03 (mmio_insufficient_data_err)
  logic          set_tx_mwr_data_payload_overrun_err; // set term for register 0x010 afu_intf_error bit(s) 02:02 (tx_mwr_data_payload_overrun_err)
  logic          set_tx_mwr_insufficient_data_err; // set term for register 0x010 afu_intf_error bit(s) 01:01 (tx_mwr_insufficient_data_err)
  logic  [10:00] vf_num_ferr_load_data; // load data for register 0x018 afu_intf_first_error bit(s) 28:18 (vf_num_ferr)
  logic  [31:00] addr_timeout_csr_reg_load_data; // load data for register 0x020 mmio_timeout_addr bit(s) 31:00 (mmio_timeout_addr)
  logic          timeout_regs_frozen_load_data; // load data for register 0x028 mmio_timeout_info bit(s) 63:63 (timeout_regs_frozen)
  logic  [07:00] tag_timeout_csr_reg_load_data; // load data for register 0x028 mmio_timeout_info bit(s) 35:28 (mmio_timeout_tag)
  logic  [09:00] dw0_len_timeout_csr_reg_load_data; // load data for register 0x028 mmio_timeout_info bit(s) 25:16 (mmio_timeout_dw0_len)
  logic  [15:00] requester_id_timeout_csr_reg_load_data; // load data for register 0x028 mmio_timeout_info bit(s) 15:00 (mmio_timeout_requester_id)
   // ******************************************************
   // *default reset value wires..
   // ******************************************************
  logic   [03:00] feature_type_default = 4'h3;
  logic           eol_default = 1'b1;
  logic   [23:00] next_dfh_byte_offset_default = 24'h0;
  logic   [03:00] feature_rev_default = 4'h2;
  logic   [11:00] feature_id_default = 12'h10;
  logic   [63:00] scratchpad_default = 64'h0;
  logic           blocking_traffic_default = 1'b0;
  logic   [10:00] vf_num_default = 11'h0;
  logic           vf_flr_access_default = 1'b0;
  logic           malformed_tlp_err_default = 1'b0;
  logic           max_payload_err_default = 1'b0;
  logic           max_read_req_size_err_default = 1'b0;
  logic           max_tag_err_default = 1'b0;
  logic           unexp_mmio_rsp_err_default = 1'b0;
  logic           mmio_timeout_err_default = 1'b0;
  logic           mmio_data_payload_overrun_err_default = 1'b0;
  logic           mmio_insufficient_data_err_default = 1'b0;
  logic           tx_mwr_data_payload_overrun_err_default = 1'b0;
  logic           tx_mwr_insufficient_data_err_default = 1'b0;
  logic   [10:00] vf_num_ferr_default = 11'h0;
  logic           vf_flr_access_ferr_default = 1'b0;
  logic           malformed_tlp_ferr_default = 1'b0;
  logic           max_payload_ferr_default = 1'b0;
  logic           max_read_req_size_ferr_default = 1'b0;
  logic           max_tag_ferr_default = 1'b0;
  logic           unexp_mmio_rsp_ferr_default = 1'b0;
  logic           mmio_timeout_ferr_default = 1'b0;
  logic           mmio_data_payload_overrun_ferr_default = 1'b0;
  logic           mmio_insufficient_data_ferr_default = 1'b0;
  logic           tx_mwr_data_payload_overrun_ferr_default = 1'b0;
  logic           tx_mwr_insufficient_data_ferr_default = 1'b0;
  logic   [31:00] mmio_timeout_addr_default = 32'h0;
  logic           timeout_regs_frozen_default = 1'b0;
  logic   [07:00] mmio_timeout_tag_default = 8'h0;
  logic   [09:00] mmio_timeout_dw0_len_default = 10'h0;
  logic   [15:00] mmio_timeout_requester_id_default = 16'h0;
  logic           tx_hdr_is_pu_mode_default = 1'b0;
  logic           mmio_immediate_frozen_default = 1'b0;
  logic   [63:00] tx_header_error_255_192_default = 64'h0;
  logic   [63:00] tx_header_error_191_128_default = 64'h0;
  logic   [63:00] tx_header_error_127_64_default = 64'h0;
  logic   [63:00] tx_header_error_63_00_default = 64'h0;
   
   // ***************************************
   // Start Manual reg and wire decls (string key for mk_cfg_module_64.pl)
   // ***************************************
   logic [7:0]      byte_en_r3;
   csr_access_type_t       csr_write_type;
   csr_access_type_t       csr_write_type_r1;
   csr_access_type_t       csr_write_type_r2;
   
   logic [HI_ADDR_BIT:02] csr_addr_r1;
   logic [07:02]          csr_addr_r2;
   logic                  csr_write_r1;
   logic                  csr_write_r2;
   logic                  core_reg_we_r3;
   logic [63:0]           csr_regwr_data_r1;
   logic [63:0]           csr_regwr_data_r2;
   logic [63:0]           csr_regwr_data_r3;
   
   logic                  csr_read_r1;
   logic                  csr_read_r2;
   logic                  csr_read_done_pulse_r2;
   logic                  csr_read_done_pulse_r3;
   logic                  csr_read_done_pulse_r4;
   
   // ######################################################################################
   // ### The wire below (rd_or_wr_r1) is a pulse used by the mk_cfg_module_64.pl script ###
   // ######################################################################################
   logic                  rd_or_wr_r1;
   
   //-------------------------------------
   // Signals
   //-------------------------------------
   ofs_fim_axi_mmio_if     csr_if();
   
   logic [HI_ADDR_BIT:0]  csr_waddr;
   logic [63:0]           csr_wdata;
   logic                  csr_write;
   
   logic [HI_ADDR_BIT:0]  csr_raddr;
   logic                  csr_read;
   logic                  csr_read_32b;
   
   // #######################################################################
   // ### The following wire names are hardcoaded into the                ###
   // ### mk_cfg_module_64.pl and is used to place the final readdata on. ###
   // #######################################################################
   logic [63:0]           csr_readdata;
   logic                  csr_readdata_valid;
   
   // #################################################################
   // ### Below here is specific to the protocol checker CSRs only. ###
   // ### It is not part of the common template                     ###
   // #################################################################
   t_prtcl_chkr_err_vector error_vector_csr;
   
   logic                  freeze_first_err_regs;
   logic                  timeout_info_regs_locked_down;
   
   // blocking traffic as a result of the protocol error logic detecting an
   // error. We never actually set this bit to one in the rtl, It is done by
   // a completion timeout that retuens all F's (signifying that we are
   // blocking traffic). The bit is only here so that is is not mistakenly
   
   // ***************************************
   // Start Manual RTL Coading (common to all templates)
   // ***************************************
   

   axi_lite2mmio axi_lite2mmio
     (
      .clk    (clk_csr),
      .rst_n  (rst_n_csr),
      .lite_if(csr_lite_if),
      .mmio_if(csr_if)
      );

   //---------------------------------
   // Map AXI write/read request to CSR write/read,
   // and send the write/read response back
   //---------------------------------
   ofs_fim_axi_csr_slave #(
      .ADDR_WIDTH ($bits(csr_waddr))
   ) mc_csr_slave (
      .csr_if             (csr_if),
      
      .csr_write          (csr_write),
      .csr_waddr          (csr_waddr),
      .csr_write_type     (csr_write_type),
      .csr_wdata          (csr_wdata),
      .csr_wstrb          (),
      
      .csr_read           (csr_read),
      .csr_raddr          (csr_raddr),
      .csr_read_32b       (csr_read_32b),
      .csr_readdata       (csr_readdata),
      .csr_readdata_valid (csr_readdata_valid)
      );
   
   always @(posedge clk_csr) begin
      csr_addr_r1             <= (csr_read ? csr_raddr[HI_ADDR_BIT:2] : csr_write ? csr_waddr[HI_ADDR_BIT:2] : csr_addr_r1); // csr_addr_r1 used my mk_cfg_module_64.pl
      csr_addr_r2             <= csr_addr_r1[07:02]; // csr_addr_r2 used my mk_cfg_module_64.pl 
      csr_write_r1            <= csr_write & rst_n_csr;
      csr_write_r2            <= csr_write_r1;
      core_reg_we_r3          <= csr_write_r2; // high fanout net Keep simple for quartus replication.
      csr_regwr_data_r1       <= csr_wdata;
      csr_regwr_data_r2       <= csr_regwr_data_r1;
      csr_regwr_data_r3       <= csr_regwr_data_r2;
      csr_read_r1             <= csr_read & ~csr_readdata_valid;
      csr_read_r2             <= csr_read_r1;
      csr_read_done_pulse_r2  <= csr_read_r1 & ~csr_read_r2;
      csr_read_done_pulse_r3  <= csr_read_done_pulse_r2;
      csr_read_done_pulse_r4  <= csr_read_done_pulse_r3;
      csr_readdata_valid      <= csr_read_done_pulse_r4;
      
      csr_write_type_r1       <= csr_write_type;
      csr_write_type_r2       <= csr_write_type_r1;
      
      
      if (csr_write_type_r2 == ofs_csr_pkg::UPPER32) begin
         byte_en_r3 <= 8'hF0;
      end else if (csr_write_type_r2 == ofs_csr_pkg::LOWER32) begin
         byte_en_r3 <= 8'h0F;
      end else if (csr_write_type_r2 == ofs_csr_pkg::FULL64) begin
         byte_en_r3 <= 8'hFF;
      end else begin
         byte_en_r3 <= 8'h00;
      end
   end // always @ (posedge clk_csr)
   
   // ######################################################################################
   // ### The wire below (rd_or_wr_r1) is a pulse used by the mk_cfg_module_64.pl script ###
   // ######################################################################################
   assign rd_or_wr_r1 = csr_read_r1 & ~csr_read_r2
                      | csr_write_r1 & ~csr_write_r2;
   
   
   // #################################################################
   // ### Below here is specific to the protocol checker CSRs only. ###
   // ### It is not part of the common template                     ###
   // #################################################################
   logic err_dcfifo_wrreq;
   logic err_dcfifo_rdreq;
   logic err_dcfifo_rdempty;

   assign err_dcfifo_wrreq = |i_error_vector;
   assign err_dcfifo_rdreq = ~err_dcfifo_rdempty;

   fim_dcfifo #(
      .DATA_WIDTH               ($bits(i_error_vector)),
      .ALMOST_FULL_THRESHOLD    (4),
      .DEPTH_RADIX              (3),
      .OVERFLOW_CHECKING_PARAM  ("OFF"),    
      .UNDERFLOW_CHECKING_PARAM ("OFF"),
      .LPM_SHOWAHEAD_PARAM      ("ON")
   ) fim_dcfifo_inst (
      .aclr      (~rst_n_csr),
      .wrclk     (clk),
      .wrreq     (|i_error_vector),
      .data      (i_error_vector),
      .wrempty   (),
      .wrfull    (),
      .wralmfull (),
      .wrusedw   (),

      .q         (error_vector_csr),
      .rdempty   (err_dcfifo_rdempty),
      .rdfull    (),
      .rdusedw   (),
      .rdclk     (clk_csr),
      .rdreq     (err_dcfifo_rdreq)
    
   );
   
   //error_vector_csr.set_tx_req_counter_oflow_err = 1'b0;                                      // 15
   assign   set_malformed_tlp_err               = error_vector_csr.malformed_tlp;               // 14
   assign   set_max_payload_err                 = error_vector_csr.max_payload;                 // 13
   assign   set_max_read_req_size_err           = error_vector_csr.max_read_req_size;           // 12
   assign   set_max_tag_err                     = error_vector_csr.max_tag;                     // 11
   //error_vector_csr.set_unaligned_addr_err    = 1'b0;                                         // 10
   //error_vector_csr.set_tag_occupied_err      = 1'b0;                                         // 09
   assign   set_unexp_mmio_rsp_err              = error_vector_csr.unexp_mmio_rsp;              // 08
   assign   set_mmio_timeout_err                = error_vector_csr.mmio_timeout;                // 07
   //error_vector_csr.set_mmio_wr_while_rst_err = 1'b0;                                         // 06
   //error_vector_csr.set_mmio_rd_while_rst_err = 1'b0;                                         // 05
   assign   set_mmio_data_payload_overrun_err   = error_vector_csr.mmio_data_payload_overrun;   // 04
   assign   set_mmio_insufficient_data_err      = error_vector_csr.mmio_insufficient_data;      // 03
   assign   set_tx_mwr_data_payload_overrun_err = error_vector_csr.tx_mwr_data_payload_overrun; // 02
   assign   set_tx_mwr_insufficient_data_err    = error_vector_csr.tx_mwr_insufficient_data;    // 01
   //error_vector_csr.set_tx_valid_violation_err    = 1'b0;                                     // 00                
   
   //----------------------------------------------------------------------------
   // FIRST ERROR signals
   //----------------------------------------------------------------------------
   assign freeze_first_err_regs = malformed_tlp_err_reg |
                                  max_payload_err_reg |
                                  max_read_req_size_err_reg |
                                  max_tag_err_reg |
                                  unexp_mmio_rsp_err_reg |
                                  mmio_timeout_err_reg |
                                  mmio_data_payload_overrun_err_reg |
                                  mmio_insufficient_data_err_reg |
                                  tx_mwr_data_payload_overrun_err_reg |
                                  tx_mwr_insufficient_data_err_reg;
   assign o_clear_errors = 0;
   
   assign vf_num_ferr_load_data = i_vf_num_load_data;
   
   assign timeout_regs_frozen_load_data = i_error_vector.mmio_timeout | timeout_info_regs_locked_down;
   
   always @(posedge clk) begin
      if (~pwr_good_clk_n) begin
         timeout_info_regs_locked_down                <= 1'b0;
      end else if (i_error_vector.mmio_timeout) begin
         timeout_info_regs_locked_down                <= 1'b1;
      end
   end

   always @(posedge clk) begin
      if (~timeout_regs_frozen_load_data) begin
         addr_timeout_csr_reg_load_data             <= i_mmio_timeout_info.addr;
         tag_timeout_csr_reg_load_data              <= i_mmio_timeout_info.tag;
         dw0_len_timeout_csr_reg_load_data          <= i_mmio_timeout_info.dw0_len;
         requester_id_timeout_csr_reg_load_data     <= i_mmio_timeout_info.requester_id;
      end
      
   end
   
   
   // BELOW IS A KEY PHRASE THE mk_cfg_module_64.pl
   // KEYS ON. DO NOT DELETE.
   // ***************************************
   // Start Auto generated rtl code
   // ***************************************
   always @(posedge clk_csr) begin
      rd_or_wr_r2 <= rd_or_wr_r1;
   end
   always @(posedge clk_csr) begin
      decode_11_8_00 <= rd_or_wr_r1 & (csr_addr_r1[11:08] == 4'h00);
      decode_11_8_01 <= rd_or_wr_r1 & (csr_addr_r1[11:08] == 4'h01);
      decode_11_8_02 <= rd_or_wr_r1 & (csr_addr_r1[11:08] == 4'h02);
      decode_11_8_03 <= rd_or_wr_r1 & (csr_addr_r1[11:08] == 4'h03);
      decode_11_8_04 <= rd_or_wr_r1 & (csr_addr_r1[11:08] == 4'h04);
      decode_11_8_05 <= rd_or_wr_r1 & (csr_addr_r1[11:08] == 4'h05);
      decode_11_8_06 <= rd_or_wr_r1 & (csr_addr_r1[11:08] == 4'h06);
      decode_11_8_07 <= rd_or_wr_r1 & (csr_addr_r1[11:08] == 4'h07);
      decode_11_8_08 <= rd_or_wr_r1 & (csr_addr_r1[11:08] == 4'h08);
      decode_11_8_09 <= rd_or_wr_r1 & (csr_addr_r1[11:08] == 4'h09);
      decode_11_8_10 <= rd_or_wr_r1 & (csr_addr_r1[11:08] == 4'h0A);
      decode_11_8_11 <= rd_or_wr_r1 & (csr_addr_r1[11:08] == 4'h0B);
      decode_11_8_12 <= rd_or_wr_r1 & (csr_addr_r1[11:08] == 4'h0C);
      decode_11_8_13 <= rd_or_wr_r1 & (csr_addr_r1[11:08] == 4'h0D);
      decode_11_8_14 <= rd_or_wr_r1 & (csr_addr_r1[11:08] == 4'h0E);
      decode_11_8_15 <= rd_or_wr_r1 & (csr_addr_r1[11:08] == 4'h0F);
   end

// *****************************************************
// RTL for the 5 bit "register" decode.
// *****************************************************
  always @(posedge clk_csr) begin
      afu_intf_dfh_en_r3                  <= rd_or_wr_r2 & decode_11_8_00 & (csr_addr_r2[07:03] == 5'b00000); // Decode for register 0x000
      afu_intf_scratchpad_en_r3           <= rd_or_wr_r2 & decode_11_8_00 & (csr_addr_r2[07:03] == 5'b00001); // Decode for register 0x008
      afu_intf_error_en_r3                <= rd_or_wr_r2 & decode_11_8_00 & (csr_addr_r2[07:03] == 5'b00010); // Decode for register 0x010
      afu_intf_first_error_en_r3          <= rd_or_wr_r2 & decode_11_8_00 & (csr_addr_r2[07:03] == 5'b00011); // Decode for register 0x018
      mmio_timeout_addr_en_r3             <= rd_or_wr_r2 & decode_11_8_00 & (csr_addr_r2[07:03] == 5'b00100); // Decode for register 0x020
      mmio_timeout_info_en_r3             <= rd_or_wr_r2 & decode_11_8_00 & (csr_addr_r2[07:03] == 5'b00101); // Decode for register 0x028
      mmio_immediate_frozen_reg_en_r3     <= rd_or_wr_r2 & decode_11_8_00 & (csr_addr_r2[07:03] == 5'b00110); // Decode for register 0x030
      mmio_tx_header_error_255_192_en_r3  <= rd_or_wr_r2 & decode_11_8_00 & (csr_addr_r2[07:03] == 5'b00111); // Decode for register 0x038
      mmio_tx_header_error_191_128_en_r3  <= rd_or_wr_r2 & decode_11_8_00 & (csr_addr_r2[07:03] == 5'b01000); // Decode for register 0x040
      mmio_tx_header_error_127_64_en_r3   <= rd_or_wr_r2 & decode_11_8_00 & (csr_addr_r2[07:03] == 5'b01001); // Decode for register 0x048
      mmio_tx_header_error_63_00_en_r3    <= rd_or_wr_r2 & decode_11_8_00 & (csr_addr_r2[07:03] == 5'b01010); // Decode for register 0x050
   end

// *****************************************************
// Start RTL for each bit and assign the 64 bit wire
// *****************************************************
// ******************************************************
// Register 0x000 afu_intf_dfh
// ******************************************************
// ******************************************************
// Bit(s) 63:60 (feature_type) of Register 0x000 afu_intf_dfh
// ******************************************************
assign feature_type_reg[03:00] = feature_type_default[03:00];
// ******************************************************
// Bit(s) 40:40 (eol) of Register 0x000 afu_intf_dfh
// ******************************************************
assign eol_reg = eol_default;
// ******************************************************
// Bit(s) 39:16 (next_dfh_byte_offset) of Register 0x000 afu_intf_dfh
// ******************************************************
assign next_dfh_byte_offset_reg[23:16] = next_dfh_byte_offset_default[23:16];
// ******************************************************
// Bit(s) 39:16 (next_dfh_byte_offset) of Register 0x000 afu_intf_dfh
// ******************************************************
assign next_dfh_byte_offset_reg[15:08] = next_dfh_byte_offset_default[15:08];
// ******************************************************
// Bit(s) 39:16 (next_dfh_byte_offset) of Register 0x000 afu_intf_dfh
// ******************************************************
assign next_dfh_byte_offset_reg[07:00] = next_dfh_byte_offset_default[07:00];
// ******************************************************
// Bit(s) 15:12 (feature_rev) of Register 0x000 afu_intf_dfh
// ******************************************************
assign feature_rev_reg[03:00] = feature_rev_default[03:00];
// ******************************************************
// Bit(s) 11:00 (feature_id) of Register 0x000 afu_intf_dfh
// ******************************************************
assign feature_id_reg[11:08] = feature_id_default[11:08];
// ******************************************************
// Bit(s) 11:00 (feature_id) of Register 0x000 afu_intf_dfh
// ******************************************************
assign feature_id_reg[07:00] = feature_id_default[07:00];

// *****************************************************
// assign the register net to all the bits.
// *****************************************************
assign afu_intf_dfh_wire = {
  feature_type_reg[03]               , feature_type_reg[02]               , feature_type_reg[01]               , feature_type_reg[00]               
, 1'b0                               , 1'b0                               , 1'b0                               , 1'b0                               
, 1'b0                               , 1'b0                               , 1'b0                               , 1'b0                               
, 1'b0                               , 1'b0                               , 1'b0                               , 1'b0                               
, 1'b0                               , 1'b0                               , 1'b0                               , 1'b0                               
, 1'b0                               , 1'b0                               , 1'b0                               , eol_reg                            
, next_dfh_byte_offset_reg[23]       , next_dfh_byte_offset_reg[22]       , next_dfh_byte_offset_reg[21]       , next_dfh_byte_offset_reg[20]       
, next_dfh_byte_offset_reg[19]       , next_dfh_byte_offset_reg[18]       , next_dfh_byte_offset_reg[17]       , next_dfh_byte_offset_reg[16]       
, next_dfh_byte_offset_reg[15]       , next_dfh_byte_offset_reg[14]       , next_dfh_byte_offset_reg[13]       , next_dfh_byte_offset_reg[12]       
, next_dfh_byte_offset_reg[11]       , next_dfh_byte_offset_reg[10]       , next_dfh_byte_offset_reg[09]       , next_dfh_byte_offset_reg[08]       
, next_dfh_byte_offset_reg[07]       , next_dfh_byte_offset_reg[06]       , next_dfh_byte_offset_reg[05]       , next_dfh_byte_offset_reg[04]       
, next_dfh_byte_offset_reg[03]       , next_dfh_byte_offset_reg[02]       , next_dfh_byte_offset_reg[01]       , next_dfh_byte_offset_reg[00]       
, feature_rev_reg[03]                , feature_rev_reg[02]                , feature_rev_reg[01]                , feature_rev_reg[00]                
, feature_id_reg[11]                 , feature_id_reg[10]                 , feature_id_reg[09]                 , feature_id_reg[08]                 
, feature_id_reg[07]                 , feature_id_reg[06]                 , feature_id_reg[05]                 , feature_id_reg[04]                 
, feature_id_reg[03]                 , feature_id_reg[02]                 , feature_id_reg[01]                 , feature_id_reg[00]                 };

// ******************************************************
// Register 0x008 afu_intf_scratchpad
// ******************************************************
// ******************************************************
// Bit(s) 63:00 (scratchpad) of Register 0x008 afu_intf_scratchpad
// ******************************************************
   always @(posedge clk_csr) begin
      if (~rst_n_csr) begin
         scratchpad_reg[63:56] <= scratchpad_default[63:56];
      end
      else if (afu_intf_scratchpad_en_r3 & core_reg_we_r3 & byte_en_r3[7]) begin
         scratchpad_reg[63:56] <= csr_regwr_data_r3[63:56];
      end
   end

// ******************************************************
// Bit(s) 63:00 (scratchpad) of Register 0x008 afu_intf_scratchpad
// ******************************************************
   always @(posedge clk_csr) begin
      if (~rst_n_csr) begin
         scratchpad_reg[55:48] <= scratchpad_default[55:48];
      end
      else if (afu_intf_scratchpad_en_r3 & core_reg_we_r3 & byte_en_r3[6]) begin
         scratchpad_reg[55:48] <= csr_regwr_data_r3[55:48];
      end
   end

// ******************************************************
// Bit(s) 63:00 (scratchpad) of Register 0x008 afu_intf_scratchpad
// ******************************************************
   always @(posedge clk_csr) begin
      if (~rst_n_csr) begin
         scratchpad_reg[47:40] <= scratchpad_default[47:40];
      end
      else if (afu_intf_scratchpad_en_r3 & core_reg_we_r3 & byte_en_r3[5]) begin
         scratchpad_reg[47:40] <= csr_regwr_data_r3[47:40];
      end
   end

// ******************************************************
// Bit(s) 63:00 (scratchpad) of Register 0x008 afu_intf_scratchpad
// ******************************************************
   always @(posedge clk_csr) begin
      if (~rst_n_csr) begin
         scratchpad_reg[39:32] <= scratchpad_default[39:32];
      end
      else if (afu_intf_scratchpad_en_r3 & core_reg_we_r3 & byte_en_r3[4]) begin
         scratchpad_reg[39:32] <= csr_regwr_data_r3[39:32];
      end
   end

// ******************************************************
// Bit(s) 63:00 (scratchpad) of Register 0x008 afu_intf_scratchpad
// ******************************************************
   always @(posedge clk_csr) begin
      if (~rst_n_csr) begin
         scratchpad_reg[31:24] <= scratchpad_default[31:24];
      end
      else if (afu_intf_scratchpad_en_r3 & core_reg_we_r3 & byte_en_r3[3]) begin
         scratchpad_reg[31:24] <= csr_regwr_data_r3[31:24];
      end
   end

// ******************************************************
// Bit(s) 63:00 (scratchpad) of Register 0x008 afu_intf_scratchpad
// ******************************************************
   always @(posedge clk_csr) begin
      if (~rst_n_csr) begin
         scratchpad_reg[23:16] <= scratchpad_default[23:16];
      end
      else if (afu_intf_scratchpad_en_r3 & core_reg_we_r3 & byte_en_r3[2]) begin
         scratchpad_reg[23:16] <= csr_regwr_data_r3[23:16];
      end
   end

// ******************************************************
// Bit(s) 63:00 (scratchpad) of Register 0x008 afu_intf_scratchpad
// ******************************************************
   always @(posedge clk_csr) begin
      if (~rst_n_csr) begin
         scratchpad_reg[15:08] <= scratchpad_default[15:08];
      end
      else if (afu_intf_scratchpad_en_r3 & core_reg_we_r3 & byte_en_r3[1]) begin
         scratchpad_reg[15:08] <= csr_regwr_data_r3[15:08];
      end
   end

// ******************************************************
// Bit(s) 63:00 (scratchpad) of Register 0x008 afu_intf_scratchpad
// ******************************************************
   always @(posedge clk_csr) begin
      if (~rst_n_csr) begin
         scratchpad_reg[07:00] <= scratchpad_default[07:00];
      end
      else if (afu_intf_scratchpad_en_r3 & core_reg_we_r3 & byte_en_r3[0]) begin
         scratchpad_reg[07:00] <= csr_regwr_data_r3[07:00];
      end
   end


// *****************************************************
// assign the register net to all the bits.
// *****************************************************
assign afu_intf_scratchpad_wire = {
  scratchpad_reg[63]                 , scratchpad_reg[62]                 , scratchpad_reg[61]                 , scratchpad_reg[60]                 
, scratchpad_reg[59]                 , scratchpad_reg[58]                 , scratchpad_reg[57]                 , scratchpad_reg[56]                 
, scratchpad_reg[55]                 , scratchpad_reg[54]                 , scratchpad_reg[53]                 , scratchpad_reg[52]                 
, scratchpad_reg[51]                 , scratchpad_reg[50]                 , scratchpad_reg[49]                 , scratchpad_reg[48]                 
, scratchpad_reg[47]                 , scratchpad_reg[46]                 , scratchpad_reg[45]                 , scratchpad_reg[44]                 
, scratchpad_reg[43]                 , scratchpad_reg[42]                 , scratchpad_reg[41]                 , scratchpad_reg[40]                 
, scratchpad_reg[39]                 , scratchpad_reg[38]                 , scratchpad_reg[37]                 , scratchpad_reg[36]                 
, scratchpad_reg[35]                 , scratchpad_reg[34]                 , scratchpad_reg[33]                 , scratchpad_reg[32]                 
, scratchpad_reg[31]                 , scratchpad_reg[30]                 , scratchpad_reg[29]                 , scratchpad_reg[28]                 
, scratchpad_reg[27]                 , scratchpad_reg[26]                 , scratchpad_reg[25]                 , scratchpad_reg[24]                 
, scratchpad_reg[23]                 , scratchpad_reg[22]                 , scratchpad_reg[21]                 , scratchpad_reg[20]                 
, scratchpad_reg[19]                 , scratchpad_reg[18]                 , scratchpad_reg[17]                 , scratchpad_reg[16]                 
, scratchpad_reg[15]                 , scratchpad_reg[14]                 , scratchpad_reg[13]                 , scratchpad_reg[12]                 
, scratchpad_reg[11]                 , scratchpad_reg[10]                 , scratchpad_reg[09]                 , scratchpad_reg[08]                 
, scratchpad_reg[07]                 , scratchpad_reg[06]                 , scratchpad_reg[05]                 , scratchpad_reg[04]                 
, scratchpad_reg[03]                 , scratchpad_reg[02]                 , scratchpad_reg[01]                 , scratchpad_reg[00]                 };

// ******************************************************
// Register 0x010 afu_intf_error
// ******************************************************
// ******************************************************
// Bit(s) 31:31 (blocking_traffic) of Register 0x010 afu_intf_error
// ******************************************************
assign blocking_traffic_reg = blocking_traffic_default;
// ******************************************************
// Bit(s) 28:18 (vf_num) of Register 0x010 afu_intf_error
// ******************************************************
   always @(posedge clk_csr) begin
      if (~rst_n_csr) begin
         vf_num_reg[10:06] <= vf_num_default[10:06];
      end
     else if (1'b1) begin
         vf_num_reg[10:06] <= i_vf_num_load_data[10:06];
       end
   end

// ******************************************************
// Bit(s) 28:18 (vf_num) of Register 0x010 afu_intf_error
// ******************************************************
   always @(posedge clk_csr) begin
      if (~rst_n_csr) begin
         vf_num_reg[05:00] <= vf_num_default[05:00];
      end
     else if (1'b1) begin
         vf_num_reg[05:00] <= i_vf_num_load_data[05:00];
       end
   end

// ******************************************************
// Bit(s) 17:17 (vf_flr_access) of Register 0x010 afu_intf_error
// ******************************************************
assign vf_flr_access_reg = vf_flr_access_default;
// ******************************************************
// Bit(s) 14:14 (malformed_tlp_err) of Register 0x010 afu_intf_error
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         malformed_tlp_err_reg <= malformed_tlp_err_default;
      end
     else if ( csr_regwr_data_r3[14] & byte_en_r3[1] & afu_intf_error_en_r3 & core_reg_we_r3) begin
         malformed_tlp_err_reg <= 1'b0;
       end
     else if (set_malformed_tlp_err) begin
         malformed_tlp_err_reg <= {1{1'b1}};
       end
   end

// ******************************************************
// Bit(s) 13:13 (max_payload_err) of Register 0x010 afu_intf_error
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         max_payload_err_reg <= max_payload_err_default;
      end
     else if ( csr_regwr_data_r3[13] & byte_en_r3[1] & afu_intf_error_en_r3 & core_reg_we_r3) begin
         max_payload_err_reg <= 1'b0;
       end
     else if (set_max_payload_err) begin
         max_payload_err_reg <= {1{1'b1}};
       end
   end

// ******************************************************
// Bit(s) 12:12 (max_read_req_size_err) of Register 0x010 afu_intf_error
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         max_read_req_size_err_reg <= max_read_req_size_err_default;
      end
     else if ( csr_regwr_data_r3[12] & byte_en_r3[1] & afu_intf_error_en_r3 & core_reg_we_r3) begin
         max_read_req_size_err_reg <= 1'b0;
       end
     else if (set_max_read_req_size_err) begin
         max_read_req_size_err_reg <= {1{1'b1}};
       end
   end

// ******************************************************
// Bit(s) 11:11 (max_tag_err) of Register 0x010 afu_intf_error
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         max_tag_err_reg <= max_tag_err_default;
      end
     else if ( csr_regwr_data_r3[11] & byte_en_r3[1] & afu_intf_error_en_r3 & core_reg_we_r3) begin
         max_tag_err_reg <= 1'b0;
       end
     else if (set_max_tag_err) begin
         max_tag_err_reg <= {1{1'b1}};
       end
   end

// ******************************************************
// Bit(s) 08:08 (unexp_mmio_rsp_err) of Register 0x010 afu_intf_error
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         unexp_mmio_rsp_err_reg <= unexp_mmio_rsp_err_default;
      end
     else if ( csr_regwr_data_r3[08] & byte_en_r3[1] & afu_intf_error_en_r3 & core_reg_we_r3) begin
         unexp_mmio_rsp_err_reg <= 1'b0;
       end
     else if (set_unexp_mmio_rsp_err) begin
         unexp_mmio_rsp_err_reg <= {1{1'b1}};
       end
   end

// ******************************************************
// Bit(s) 07:07 (mmio_timeout_err) of Register 0x010 afu_intf_error
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         mmio_timeout_err_reg <= mmio_timeout_err_default;
      end
     else if ( csr_regwr_data_r3[07] & byte_en_r3[0] & afu_intf_error_en_r3 & core_reg_we_r3) begin
         mmio_timeout_err_reg <= 1'b0;
       end
     else if (set_mmio_timeout_err) begin
         mmio_timeout_err_reg <= {1{1'b1}};
       end
   end

// ******************************************************
// Bit(s) 04:04 (mmio_data_payload_overrun_err) of Register 0x010 afu_intf_error
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         mmio_data_payload_overrun_err_reg <= mmio_data_payload_overrun_err_default;
      end
     else if ( csr_regwr_data_r3[04] & byte_en_r3[0] & afu_intf_error_en_r3 & core_reg_we_r3) begin
         mmio_data_payload_overrun_err_reg <= 1'b0;
       end
     else if (set_mmio_data_payload_overrun_err) begin
         mmio_data_payload_overrun_err_reg <= {1{1'b1}};
       end
   end

// ******************************************************
// Bit(s) 03:03 (mmio_insufficient_data_err) of Register 0x010 afu_intf_error
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         mmio_insufficient_data_err_reg <= mmio_insufficient_data_err_default;
      end
     else if ( csr_regwr_data_r3[03] & byte_en_r3[0] & afu_intf_error_en_r3 & core_reg_we_r3) begin
         mmio_insufficient_data_err_reg <= 1'b0;
       end
     else if (set_mmio_insufficient_data_err) begin
         mmio_insufficient_data_err_reg <= {1{1'b1}};
       end
   end

// ******************************************************
// Bit(s) 02:02 (tx_mwr_data_payload_overrun_err) of Register 0x010 afu_intf_error
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         tx_mwr_data_payload_overrun_err_reg <= tx_mwr_data_payload_overrun_err_default;
      end
     else if ( csr_regwr_data_r3[02] & byte_en_r3[0] & afu_intf_error_en_r3 & core_reg_we_r3) begin
         tx_mwr_data_payload_overrun_err_reg <= 1'b0;
       end
     else if (set_tx_mwr_data_payload_overrun_err) begin
         tx_mwr_data_payload_overrun_err_reg <= {1{1'b1}};
       end
   end

// ******************************************************
// Bit(s) 01:01 (tx_mwr_insufficient_data_err) of Register 0x010 afu_intf_error
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         tx_mwr_insufficient_data_err_reg <= tx_mwr_insufficient_data_err_default;
      end
     else if ( csr_regwr_data_r3[01] & byte_en_r3[0] & afu_intf_error_en_r3 & core_reg_we_r3) begin
         tx_mwr_insufficient_data_err_reg <= 1'b0;
       end
     else if (set_tx_mwr_insufficient_data_err) begin
         tx_mwr_insufficient_data_err_reg <= {1{1'b1}};
       end
   end


// *****************************************************
// assign the register net to all the bits.
// *****************************************************
assign afu_intf_error_wire = {
  1'b0                               , 1'b0                               , 1'b0                               , 1'b0                               
, 1'b0                               , 1'b0                               , 1'b0                               , 1'b0                               
, 1'b0                               , 1'b0                               , 1'b0                               , 1'b0                               
, 1'b0                               , 1'b0                               , 1'b0                               , 1'b0                               
, 1'b0                               , 1'b0                               , 1'b0                               , 1'b0                               
, 1'b0                               , 1'b0                               , 1'b0                               , 1'b0                               
, 1'b0                               , 1'b0                               , 1'b0                               , 1'b0                               
, 1'b0                               , 1'b0                               , 1'b0                               , 1'b0                               
, blocking_traffic_reg               , 1'b0                               , 1'b0                               , vf_num_reg[10]                     
, vf_num_reg[09]                     , vf_num_reg[08]                     , vf_num_reg[07]                     , vf_num_reg[06]                     
, vf_num_reg[05]                     , vf_num_reg[04]                     , vf_num_reg[03]                     , vf_num_reg[02]                     
, vf_num_reg[01]                     , vf_num_reg[00]                     , vf_flr_access_reg                  , 1'b0                               
, 1'b0                               , malformed_tlp_err_reg              , max_payload_err_reg                , max_read_req_size_err_reg          
, max_tag_err_reg                    , 1'b0                               , 1'b0                               , unexp_mmio_rsp_err_reg             
, mmio_timeout_err_reg               , 1'b0                               , 1'b0                               , mmio_data_payload_overrun_err_reg  
, mmio_insufficient_data_err_reg     , tx_mwr_data_payload_overrun_err_reg, tx_mwr_insufficient_data_err_reg   , 1'b0                               };

// ******************************************************
// Register 0x018 afu_intf_first_error
// ******************************************************
// ******************************************************
// Bit(s) 28:18 (vf_num_ferr) of Register 0x018 afu_intf_first_error
// ******************************************************
   always @(posedge clk_csr) begin
      if (~rst_n_csr) begin
         vf_num_ferr_reg[10:06] <= vf_num_ferr_default[10:06];
      end
     else if (1'b1) begin
         vf_num_ferr_reg[10:06] <= vf_num_ferr_load_data[10:06];
       end
   end

// ******************************************************
// Bit(s) 28:18 (vf_num_ferr) of Register 0x018 afu_intf_first_error
// ******************************************************
   always @(posedge clk_csr) begin
      if (~rst_n_csr) begin
         vf_num_ferr_reg[05:00] <= vf_num_ferr_default[05:00];
      end
     else if (1'b1) begin
         vf_num_ferr_reg[05:00] <= vf_num_ferr_load_data[05:00];
       end
   end

// ******************************************************
// Bit(s) 17:17 (vf_flr_access_ferr) of Register 0x018 afu_intf_first_error
// ******************************************************
assign vf_flr_access_ferr_reg = vf_flr_access_ferr_default;
// ******************************************************
// Bit(s) 14:14 (malformed_tlp_ferr) of Register 0x018 afu_intf_first_error
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         malformed_tlp_ferr_reg <= malformed_tlp_ferr_default;
      end
     else if ( csr_regwr_data_r3[14] & byte_en_r3[1] & afu_intf_first_error_en_r3 & core_reg_we_r3) begin
         malformed_tlp_ferr_reg <= 1'b0;
       end
     else if (set_malformed_tlp_err & ~freeze_first_err_regs) begin
         malformed_tlp_ferr_reg <= {1{1'b1}};
       end
     else if (~set_malformed_tlp_err & ~freeze_first_err_regs) begin
         malformed_tlp_ferr_reg <= {1{1'b0}};
       end
   end

// ******************************************************
// Bit(s) 13:13 (max_payload_ferr) of Register 0x018 afu_intf_first_error
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         max_payload_ferr_reg <= max_payload_ferr_default;
      end
     else if ( csr_regwr_data_r3[13] & byte_en_r3[1] & afu_intf_first_error_en_r3 & core_reg_we_r3) begin
         max_payload_ferr_reg <= 1'b0;
       end
     else if (set_max_payload_err & ~freeze_first_err_regs) begin
         max_payload_ferr_reg <= {1{1'b1}};
       end
     else if (~set_max_payload_err & ~freeze_first_err_regs) begin
         max_payload_ferr_reg <= {1{1'b0}};
       end
   end

// ******************************************************
// Bit(s) 12:12 (max_read_req_size_ferr) of Register 0x018 afu_intf_first_error
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         max_read_req_size_ferr_reg <= max_read_req_size_ferr_default;
      end
     else if ( csr_regwr_data_r3[12] & byte_en_r3[1] & afu_intf_first_error_en_r3 & core_reg_we_r3) begin
         max_read_req_size_ferr_reg <= 1'b0;
       end
     else if (set_max_read_req_size_err & ~freeze_first_err_regs) begin
         max_read_req_size_ferr_reg <= {1{1'b1}};
       end
     else if (~set_max_read_req_size_err & ~freeze_first_err_regs) begin
         max_read_req_size_ferr_reg <= {1{1'b0}};
       end
   end

// ******************************************************
// Bit(s) 11:11 (max_tag_ferr) of Register 0x018 afu_intf_first_error
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         max_tag_ferr_reg <= max_tag_ferr_default;
      end
     else if ( csr_regwr_data_r3[11] & byte_en_r3[1] & afu_intf_first_error_en_r3 & core_reg_we_r3) begin
         max_tag_ferr_reg <= 1'b0;
       end
     else if (set_max_tag_err & ~freeze_first_err_regs) begin
         max_tag_ferr_reg <= {1{1'b1}};
       end
     else if (~set_max_tag_err & ~freeze_first_err_regs) begin
         max_tag_ferr_reg <= {1{1'b0}};
       end
   end

// ******************************************************
// Bit(s) 08:08 (unexp_mmio_rsp_ferr) of Register 0x018 afu_intf_first_error
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         unexp_mmio_rsp_ferr_reg <= unexp_mmio_rsp_ferr_default;
      end
     else if ( csr_regwr_data_r3[08] & byte_en_r3[1] & afu_intf_first_error_en_r3 & core_reg_we_r3) begin
         unexp_mmio_rsp_ferr_reg <= 1'b0;
       end
     else if (set_unexp_mmio_rsp_err & ~freeze_first_err_regs) begin
         unexp_mmio_rsp_ferr_reg <= {1{1'b1}};
       end
     else if (~set_unexp_mmio_rsp_err & ~freeze_first_err_regs) begin
         unexp_mmio_rsp_ferr_reg <= {1{1'b0}};
       end
   end

// ******************************************************
// Bit(s) 07:07 (mmio_timeout_ferr) of Register 0x018 afu_intf_first_error
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         mmio_timeout_ferr_reg <= mmio_timeout_ferr_default;
      end
     else if ( csr_regwr_data_r3[07] & byte_en_r3[0] & afu_intf_first_error_en_r3 & core_reg_we_r3) begin
         mmio_timeout_ferr_reg <= 1'b0;
       end
     else if (set_mmio_timeout_err & ~freeze_first_err_regs) begin
         mmio_timeout_ferr_reg <= {1{1'b1}};
       end
     else if (~set_mmio_timeout_err & ~freeze_first_err_regs) begin
         mmio_timeout_ferr_reg <= {1{1'b0}};
       end
   end

// ******************************************************
// Bit(s) 04:04 (mmio_data_payload_overrun_ferr) of Register 0x018 afu_intf_first_error
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         mmio_data_payload_overrun_ferr_reg <= mmio_data_payload_overrun_ferr_default;
      end
     else if ( csr_regwr_data_r3[04] & byte_en_r3[0] & afu_intf_first_error_en_r3 & core_reg_we_r3) begin
         mmio_data_payload_overrun_ferr_reg <= 1'b0;
       end
     else if (set_mmio_data_payload_overrun_err & ~freeze_first_err_regs) begin
         mmio_data_payload_overrun_ferr_reg <= {1{1'b1}};
       end
     else if (~set_mmio_data_payload_overrun_err & ~freeze_first_err_regs) begin
         mmio_data_payload_overrun_ferr_reg <= {1{1'b0}};
       end
   end

// ******************************************************
// Bit(s) 03:03 (mmio_insufficient_data_ferr) of Register 0x018 afu_intf_first_error
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         mmio_insufficient_data_ferr_reg <= mmio_insufficient_data_ferr_default;
      end
     else if ( csr_regwr_data_r3[03] & byte_en_r3[0] & afu_intf_first_error_en_r3 & core_reg_we_r3) begin
         mmio_insufficient_data_ferr_reg <= 1'b0;
       end
     else if (set_mmio_insufficient_data_err & ~freeze_first_err_regs) begin
         mmio_insufficient_data_ferr_reg <= {1{1'b1}};
       end
     else if (~set_mmio_insufficient_data_err & ~freeze_first_err_regs) begin
         mmio_insufficient_data_ferr_reg <= {1{1'b0}};
       end
   end

// ******************************************************
// Bit(s) 02:02 (tx_mwr_data_payload_overrun_ferr) of Register 0x018 afu_intf_first_error
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         tx_mwr_data_payload_overrun_ferr_reg <= tx_mwr_data_payload_overrun_ferr_default;
      end
     else if ( csr_regwr_data_r3[02] & byte_en_r3[0] & afu_intf_first_error_en_r3 & core_reg_we_r3) begin
         tx_mwr_data_payload_overrun_ferr_reg <= 1'b0;
       end
     else if (set_tx_mwr_data_payload_overrun_err & ~freeze_first_err_regs) begin
         tx_mwr_data_payload_overrun_ferr_reg <= {1{1'b1}};
       end
     else if (~set_tx_mwr_data_payload_overrun_err & ~freeze_first_err_regs) begin
         tx_mwr_data_payload_overrun_ferr_reg <= {1{1'b0}};
       end
   end

// ******************************************************
// Bit(s) 01:01 (tx_mwr_insufficient_data_ferr) of Register 0x018 afu_intf_first_error
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         tx_mwr_insufficient_data_ferr_reg <= tx_mwr_insufficient_data_ferr_default;
      end
     else if ( csr_regwr_data_r3[01] & byte_en_r3[0] & afu_intf_first_error_en_r3 & core_reg_we_r3) begin
         tx_mwr_insufficient_data_ferr_reg <= 1'b0;
       end
     else if (set_tx_mwr_insufficient_data_err & ~freeze_first_err_regs) begin
         tx_mwr_insufficient_data_ferr_reg <= {1{1'b1}};
       end
     else if (~set_tx_mwr_insufficient_data_err & ~freeze_first_err_regs) begin
         tx_mwr_insufficient_data_ferr_reg <= {1{1'b0}};
       end
   end


// *****************************************************
// assign the register net to all the bits.
// *****************************************************
assign afu_intf_first_error_wire = {
  1'b0                               , 1'b0                               , 1'b0                               , 1'b0                               
, 1'b0                               , 1'b0                               , 1'b0                               , 1'b0                               
, 1'b0                               , 1'b0                               , 1'b0                               , 1'b0                               
, 1'b0                               , 1'b0                               , 1'b0                               , 1'b0                               
, 1'b0                               , 1'b0                               , 1'b0                               , 1'b0                               
, 1'b0                               , 1'b0                               , 1'b0                               , 1'b0                               
, 1'b0                               , 1'b0                               , 1'b0                               , 1'b0                               
, 1'b0                               , 1'b0                               , 1'b0                               , 1'b0                               
, 1'b0                               , 1'b0                               , 1'b0                               , vf_num_ferr_reg[10]                
, vf_num_ferr_reg[09]                , vf_num_ferr_reg[08]                , vf_num_ferr_reg[07]                , vf_num_ferr_reg[06]                
, vf_num_ferr_reg[05]                , vf_num_ferr_reg[04]                , vf_num_ferr_reg[03]                , vf_num_ferr_reg[02]                
, vf_num_ferr_reg[01]                , vf_num_ferr_reg[00]                , vf_flr_access_ferr_reg             , 1'b0                               
, 1'b0                               , malformed_tlp_ferr_reg             , max_payload_ferr_reg               , max_read_req_size_ferr_reg         
, max_tag_ferr_reg                   , 1'b0                               , 1'b0                               , unexp_mmio_rsp_ferr_reg            
, mmio_timeout_ferr_reg              , 1'b0                               , 1'b0                               , mmio_data_payload_overrun_ferr_reg 
, mmio_insufficient_data_ferr_reg    , tx_mwr_data_payload_overrun_ferr_reg, tx_mwr_insufficient_data_ferr_reg  , 1'b0                               };

// ******************************************************
// Register 0x020 mmio_timeout_addr
// ******************************************************
// ******************************************************
// Bit(s) 31:00 (mmio_timeout_addr) of Register 0x020 mmio_timeout_addr
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         mmio_timeout_addr_reg[31:24] <= mmio_timeout_addr_default[31:24];
      end
     else if (1'b1) begin
         mmio_timeout_addr_reg[31:24] <= addr_timeout_csr_reg_load_data[31:24];
       end
   end

// ******************************************************
// Bit(s) 31:00 (mmio_timeout_addr) of Register 0x020 mmio_timeout_addr
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         mmio_timeout_addr_reg[23:16] <= mmio_timeout_addr_default[23:16];
      end
     else if (1'b1) begin
         mmio_timeout_addr_reg[23:16] <= addr_timeout_csr_reg_load_data[23:16];
       end
   end

// ******************************************************
// Bit(s) 31:00 (mmio_timeout_addr) of Register 0x020 mmio_timeout_addr
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         mmio_timeout_addr_reg[15:08] <= mmio_timeout_addr_default[15:08];
      end
     else if (1'b1) begin
         mmio_timeout_addr_reg[15:08] <= addr_timeout_csr_reg_load_data[15:08];
       end
   end

// ******************************************************
// Bit(s) 31:00 (mmio_timeout_addr) of Register 0x020 mmio_timeout_addr
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         mmio_timeout_addr_reg[07:00] <= mmio_timeout_addr_default[07:00];
      end
     else if (1'b1) begin
         mmio_timeout_addr_reg[07:00] <= addr_timeout_csr_reg_load_data[07:00];
       end
   end


// *****************************************************
// assign the register net to all the bits.
// *****************************************************
assign mmio_timeout_addr_wire = {
  1'b0                               , 1'b0                               , 1'b0                               , 1'b0                               
, 1'b0                               , 1'b0                               , 1'b0                               , 1'b0                               
, 1'b0                               , 1'b0                               , 1'b0                               , 1'b0                               
, 1'b0                               , 1'b0                               , 1'b0                               , 1'b0                               
, 1'b0                               , 1'b0                               , 1'b0                               , 1'b0                               
, 1'b0                               , 1'b0                               , 1'b0                               , 1'b0                               
, 1'b0                               , 1'b0                               , 1'b0                               , 1'b0                               
, 1'b0                               , 1'b0                               , 1'b0                               , 1'b0                               
, mmio_timeout_addr_reg[31]          , mmio_timeout_addr_reg[30]          , mmio_timeout_addr_reg[29]          , mmio_timeout_addr_reg[28]          
, mmio_timeout_addr_reg[27]          , mmio_timeout_addr_reg[26]          , mmio_timeout_addr_reg[25]          , mmio_timeout_addr_reg[24]          
, mmio_timeout_addr_reg[23]          , mmio_timeout_addr_reg[22]          , mmio_timeout_addr_reg[21]          , mmio_timeout_addr_reg[20]          
, mmio_timeout_addr_reg[19]          , mmio_timeout_addr_reg[18]          , mmio_timeout_addr_reg[17]          , mmio_timeout_addr_reg[16]          
, mmio_timeout_addr_reg[15]          , mmio_timeout_addr_reg[14]          , mmio_timeout_addr_reg[13]          , mmio_timeout_addr_reg[12]          
, mmio_timeout_addr_reg[11]          , mmio_timeout_addr_reg[10]          , mmio_timeout_addr_reg[09]          , mmio_timeout_addr_reg[08]          
, mmio_timeout_addr_reg[07]          , mmio_timeout_addr_reg[06]          , mmio_timeout_addr_reg[05]          , mmio_timeout_addr_reg[04]          
, mmio_timeout_addr_reg[03]          , mmio_timeout_addr_reg[02]          , mmio_timeout_addr_reg[01]          , mmio_timeout_addr_reg[00]          };

// ******************************************************
// Register 0x028 mmio_timeout_info
// ******************************************************
// ******************************************************
// Bit(s) 63:63 (timeout_regs_frozen) of Register 0x028 mmio_timeout_info
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         timeout_regs_frozen_reg <= timeout_regs_frozen_default;
      end
     else if (1'b1) begin
         timeout_regs_frozen_reg <= timeout_regs_frozen_load_data;
       end
   end

// ******************************************************
// Bit(s) 35:28 (mmio_timeout_tag) of Register 0x028 mmio_timeout_info
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         mmio_timeout_tag_reg[07:04] <= mmio_timeout_tag_default[07:04];
      end
     else if (1'b1) begin
         mmio_timeout_tag_reg[07:04] <= tag_timeout_csr_reg_load_data[07:04];
       end
   end

// ******************************************************
// Bit(s) 35:28 (mmio_timeout_tag) of Register 0x028 mmio_timeout_info
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         mmio_timeout_tag_reg[03:00] <= mmio_timeout_tag_default[03:00];
      end
     else if (1'b1) begin
         mmio_timeout_tag_reg[03:00] <= tag_timeout_csr_reg_load_data[03:00];
       end
   end

// ******************************************************
// Bit(s) 25:16 (mmio_timeout_dw0_len) of Register 0x028 mmio_timeout_info
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         mmio_timeout_dw0_len_reg[09:08] <= mmio_timeout_dw0_len_default[09:08];
      end
     else if (1'b1) begin
         mmio_timeout_dw0_len_reg[09:08] <= dw0_len_timeout_csr_reg_load_data[09:08];
       end
   end

// ******************************************************
// Bit(s) 25:16 (mmio_timeout_dw0_len) of Register 0x028 mmio_timeout_info
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         mmio_timeout_dw0_len_reg[07:00] <= mmio_timeout_dw0_len_default[07:00];
      end
     else if (1'b1) begin
         mmio_timeout_dw0_len_reg[07:00] <= dw0_len_timeout_csr_reg_load_data[07:00];
       end
   end

// ******************************************************
// Bit(s) 15:00 (mmio_timeout_requester_id) of Register 0x028 mmio_timeout_info
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         mmio_timeout_requester_id_reg[15:08] <= mmio_timeout_requester_id_default[15:08];
      end
     else if (1'b1) begin
         mmio_timeout_requester_id_reg[15:08] <= requester_id_timeout_csr_reg_load_data[15:08];
       end
   end

// ******************************************************
// Bit(s) 15:00 (mmio_timeout_requester_id) of Register 0x028 mmio_timeout_info
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         mmio_timeout_requester_id_reg[07:00] <= mmio_timeout_requester_id_default[07:00];
      end
     else if (1'b1) begin
         mmio_timeout_requester_id_reg[07:00] <= requester_id_timeout_csr_reg_load_data[07:00];
       end
   end


// *****************************************************
// assign the register net to all the bits.
// *****************************************************
assign mmio_timeout_info_wire = {
  timeout_regs_frozen_reg            , 1'b0                               , 1'b0                               , 1'b0                               
, 1'b0                               , 1'b0                               , 1'b0                               , 1'b0                               
, 1'b0                               , 1'b0                               , 1'b0                               , 1'b0                               
, 1'b0                               , 1'b0                               , 1'b0                               , 1'b0                               
, 1'b0                               , 1'b0                               , 1'b0                               , 1'b0                               
, 1'b0                               , 1'b0                               , 1'b0                               , 1'b0                               
, 1'b0                               , 1'b0                               , 1'b0                               , 1'b0                               
, mmio_timeout_tag_reg[07]           , mmio_timeout_tag_reg[06]           , mmio_timeout_tag_reg[05]           , mmio_timeout_tag_reg[04]           
, mmio_timeout_tag_reg[03]           , mmio_timeout_tag_reg[02]           , mmio_timeout_tag_reg[01]           , mmio_timeout_tag_reg[00]           
, 1'b0                               , 1'b0                               , mmio_timeout_dw0_len_reg[09]       , mmio_timeout_dw0_len_reg[08]       
, mmio_timeout_dw0_len_reg[07]       , mmio_timeout_dw0_len_reg[06]       , mmio_timeout_dw0_len_reg[05]       , mmio_timeout_dw0_len_reg[04]       
, mmio_timeout_dw0_len_reg[03]       , mmio_timeout_dw0_len_reg[02]       , mmio_timeout_dw0_len_reg[01]       , mmio_timeout_dw0_len_reg[00]       
, mmio_timeout_requester_id_reg[15]  , mmio_timeout_requester_id_reg[14]  , mmio_timeout_requester_id_reg[13]  , mmio_timeout_requester_id_reg[12]  
, mmio_timeout_requester_id_reg[11]  , mmio_timeout_requester_id_reg[10]  , mmio_timeout_requester_id_reg[09]  , mmio_timeout_requester_id_reg[08]  
, mmio_timeout_requester_id_reg[07]  , mmio_timeout_requester_id_reg[06]  , mmio_timeout_requester_id_reg[05]  , mmio_timeout_requester_id_reg[04]  
, mmio_timeout_requester_id_reg[03]  , mmio_timeout_requester_id_reg[02]  , mmio_timeout_requester_id_reg[01]  , mmio_timeout_requester_id_reg[00]  };

// ******************************************************
// Register 0x030 mmio_immediate_frozen_reg
// ******************************************************
// ******************************************************
// Bit(s) 01:01 (tx_hdr_is_pu_mode) of Register 0x030 mmio_immediate_frozen_reg
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         tx_hdr_is_pu_mode_reg <= tx_hdr_is_pu_mode_default;
      end
     else if (1'b1) begin
         tx_hdr_is_pu_mode_reg <= i_tx_hdr_is_pu_mode_load_data;
       end
   end

// ******************************************************
// Bit(s) 00:00 (mmio_immediate_frozen) of Register 0x030 mmio_immediate_frozen_reg
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         mmio_immediate_frozen_reg <= mmio_immediate_frozen_default;
      end
     else if (1'b1) begin
         mmio_immediate_frozen_reg <= i_mmio_immediate_frozen_load_data;
       end
   end


// *****************************************************
// assign the register net to all the bits.
// *****************************************************
assign mmio_immediate_frozen_reg_wire = {
  1'b0                               , 1'b0                               , 1'b0                               , 1'b0                               
, 1'b0                               , 1'b0                               , 1'b0                               , 1'b0                               
, 1'b0                               , 1'b0                               , 1'b0                               , 1'b0                               
, 1'b0                               , 1'b0                               , 1'b0                               , 1'b0                               
, 1'b0                               , 1'b0                               , 1'b0                               , 1'b0                               
, 1'b0                               , 1'b0                               , 1'b0                               , 1'b0                               
, 1'b0                               , 1'b0                               , 1'b0                               , 1'b0                               
, 1'b0                               , 1'b0                               , 1'b0                               , 1'b0                               
, 1'b0                               , 1'b0                               , 1'b0                               , 1'b0                               
, 1'b0                               , 1'b0                               , 1'b0                               , 1'b0                               
, 1'b0                               , 1'b0                               , 1'b0                               , 1'b0                               
, 1'b0                               , 1'b0                               , 1'b0                               , 1'b0                               
, 1'b0                               , 1'b0                               , 1'b0                               , 1'b0                               
, 1'b0                               , 1'b0                               , 1'b0                               , 1'b0                               
, 1'b0                               , 1'b0                               , 1'b0                               , 1'b0                               
, 1'b0                               , 1'b0                               , tx_hdr_is_pu_mode_reg              , mmio_immediate_frozen_reg          };

// ******************************************************
// Register 0x038 mmio_tx_header_error_255_192
// ******************************************************
// ******************************************************
// Bit(s) 63:00 (tx_header_error_255_192) of Register 0x038 mmio_tx_header_error_255_192
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         tx_header_error_255_192_reg[63:56] <= tx_header_error_255_192_default[63:56];
      end
     else if (1'b1) begin
         tx_header_error_255_192_reg[63:56] <= i_tx_header_error_255_192_load_data[63:56];
       end
   end

// ******************************************************
// Bit(s) 63:00 (tx_header_error_255_192) of Register 0x038 mmio_tx_header_error_255_192
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         tx_header_error_255_192_reg[55:48] <= tx_header_error_255_192_default[55:48];
      end
     else if (1'b1) begin
         tx_header_error_255_192_reg[55:48] <= i_tx_header_error_255_192_load_data[55:48];
       end
   end

// ******************************************************
// Bit(s) 63:00 (tx_header_error_255_192) of Register 0x038 mmio_tx_header_error_255_192
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         tx_header_error_255_192_reg[47:40] <= tx_header_error_255_192_default[47:40];
      end
     else if (1'b1) begin
         tx_header_error_255_192_reg[47:40] <= i_tx_header_error_255_192_load_data[47:40];
       end
   end

// ******************************************************
// Bit(s) 63:00 (tx_header_error_255_192) of Register 0x038 mmio_tx_header_error_255_192
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         tx_header_error_255_192_reg[39:32] <= tx_header_error_255_192_default[39:32];
      end
     else if (1'b1) begin
         tx_header_error_255_192_reg[39:32] <= i_tx_header_error_255_192_load_data[39:32];
       end
   end

// ******************************************************
// Bit(s) 63:00 (tx_header_error_255_192) of Register 0x038 mmio_tx_header_error_255_192
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         tx_header_error_255_192_reg[31:24] <= tx_header_error_255_192_default[31:24];
      end
     else if (1'b1) begin
         tx_header_error_255_192_reg[31:24] <= i_tx_header_error_255_192_load_data[31:24];
       end
   end

// ******************************************************
// Bit(s) 63:00 (tx_header_error_255_192) of Register 0x038 mmio_tx_header_error_255_192
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         tx_header_error_255_192_reg[23:16] <= tx_header_error_255_192_default[23:16];
      end
     else if (1'b1) begin
         tx_header_error_255_192_reg[23:16] <= i_tx_header_error_255_192_load_data[23:16];
       end
   end

// ******************************************************
// Bit(s) 63:00 (tx_header_error_255_192) of Register 0x038 mmio_tx_header_error_255_192
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         tx_header_error_255_192_reg[15:08] <= tx_header_error_255_192_default[15:08];
      end
     else if (1'b1) begin
         tx_header_error_255_192_reg[15:08] <= i_tx_header_error_255_192_load_data[15:08];
       end
   end

// ******************************************************
// Bit(s) 63:00 (tx_header_error_255_192) of Register 0x038 mmio_tx_header_error_255_192
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         tx_header_error_255_192_reg[07:00] <= tx_header_error_255_192_default[07:00];
      end
     else if (1'b1) begin
         tx_header_error_255_192_reg[07:00] <= i_tx_header_error_255_192_load_data[07:00];
       end
   end


// *****************************************************
// assign the register net to all the bits.
// *****************************************************
assign mmio_tx_header_error_255_192_wire = {
  tx_header_error_255_192_reg[63]    , tx_header_error_255_192_reg[62]    , tx_header_error_255_192_reg[61]    , tx_header_error_255_192_reg[60]    
, tx_header_error_255_192_reg[59]    , tx_header_error_255_192_reg[58]    , tx_header_error_255_192_reg[57]    , tx_header_error_255_192_reg[56]    
, tx_header_error_255_192_reg[55]    , tx_header_error_255_192_reg[54]    , tx_header_error_255_192_reg[53]    , tx_header_error_255_192_reg[52]    
, tx_header_error_255_192_reg[51]    , tx_header_error_255_192_reg[50]    , tx_header_error_255_192_reg[49]    , tx_header_error_255_192_reg[48]    
, tx_header_error_255_192_reg[47]    , tx_header_error_255_192_reg[46]    , tx_header_error_255_192_reg[45]    , tx_header_error_255_192_reg[44]    
, tx_header_error_255_192_reg[43]    , tx_header_error_255_192_reg[42]    , tx_header_error_255_192_reg[41]    , tx_header_error_255_192_reg[40]    
, tx_header_error_255_192_reg[39]    , tx_header_error_255_192_reg[38]    , tx_header_error_255_192_reg[37]    , tx_header_error_255_192_reg[36]    
, tx_header_error_255_192_reg[35]    , tx_header_error_255_192_reg[34]    , tx_header_error_255_192_reg[33]    , tx_header_error_255_192_reg[32]    
, tx_header_error_255_192_reg[31]    , tx_header_error_255_192_reg[30]    , tx_header_error_255_192_reg[29]    , tx_header_error_255_192_reg[28]    
, tx_header_error_255_192_reg[27]    , tx_header_error_255_192_reg[26]    , tx_header_error_255_192_reg[25]    , tx_header_error_255_192_reg[24]    
, tx_header_error_255_192_reg[23]    , tx_header_error_255_192_reg[22]    , tx_header_error_255_192_reg[21]    , tx_header_error_255_192_reg[20]    
, tx_header_error_255_192_reg[19]    , tx_header_error_255_192_reg[18]    , tx_header_error_255_192_reg[17]    , tx_header_error_255_192_reg[16]    
, tx_header_error_255_192_reg[15]    , tx_header_error_255_192_reg[14]    , tx_header_error_255_192_reg[13]    , tx_header_error_255_192_reg[12]    
, tx_header_error_255_192_reg[11]    , tx_header_error_255_192_reg[10]    , tx_header_error_255_192_reg[09]    , tx_header_error_255_192_reg[08]    
, tx_header_error_255_192_reg[07]    , tx_header_error_255_192_reg[06]    , tx_header_error_255_192_reg[05]    , tx_header_error_255_192_reg[04]    
, tx_header_error_255_192_reg[03]    , tx_header_error_255_192_reg[02]    , tx_header_error_255_192_reg[01]    , tx_header_error_255_192_reg[00]    };

// ******************************************************
// Register 0x040 mmio_tx_header_error_191_128
// ******************************************************
// ******************************************************
// Bit(s) 63:00 (tx_header_error_191_128) of Register 0x040 mmio_tx_header_error_191_128
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         tx_header_error_191_128_reg[63:56] <= tx_header_error_191_128_default[63:56];
      end
     else if (1'b1) begin
         tx_header_error_191_128_reg[63:56] <= i_tx_header_error_191_128_load_data[63:56];
       end
   end

// ******************************************************
// Bit(s) 63:00 (tx_header_error_191_128) of Register 0x040 mmio_tx_header_error_191_128
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         tx_header_error_191_128_reg[55:48] <= tx_header_error_191_128_default[55:48];
      end
     else if (1'b1) begin
         tx_header_error_191_128_reg[55:48] <= i_tx_header_error_191_128_load_data[55:48];
       end
   end

// ******************************************************
// Bit(s) 63:00 (tx_header_error_191_128) of Register 0x040 mmio_tx_header_error_191_128
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         tx_header_error_191_128_reg[47:40] <= tx_header_error_191_128_default[47:40];
      end
     else if (1'b1) begin
         tx_header_error_191_128_reg[47:40] <= i_tx_header_error_191_128_load_data[47:40];
       end
   end

// ******************************************************
// Bit(s) 63:00 (tx_header_error_191_128) of Register 0x040 mmio_tx_header_error_191_128
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         tx_header_error_191_128_reg[39:32] <= tx_header_error_191_128_default[39:32];
      end
     else if (1'b1) begin
         tx_header_error_191_128_reg[39:32] <= i_tx_header_error_191_128_load_data[39:32];
       end
   end

// ******************************************************
// Bit(s) 63:00 (tx_header_error_191_128) of Register 0x040 mmio_tx_header_error_191_128
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         tx_header_error_191_128_reg[31:24] <= tx_header_error_191_128_default[31:24];
      end
     else if (1'b1) begin
         tx_header_error_191_128_reg[31:24] <= i_tx_header_error_191_128_load_data[31:24];
       end
   end

// ******************************************************
// Bit(s) 63:00 (tx_header_error_191_128) of Register 0x040 mmio_tx_header_error_191_128
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         tx_header_error_191_128_reg[23:16] <= tx_header_error_191_128_default[23:16];
      end
     else if (1'b1) begin
         tx_header_error_191_128_reg[23:16] <= i_tx_header_error_191_128_load_data[23:16];
       end
   end

// ******************************************************
// Bit(s) 63:00 (tx_header_error_191_128) of Register 0x040 mmio_tx_header_error_191_128
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         tx_header_error_191_128_reg[15:08] <= tx_header_error_191_128_default[15:08];
      end
     else if (1'b1) begin
         tx_header_error_191_128_reg[15:08] <= i_tx_header_error_191_128_load_data[15:08];
       end
   end

// ******************************************************
// Bit(s) 63:00 (tx_header_error_191_128) of Register 0x040 mmio_tx_header_error_191_128
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         tx_header_error_191_128_reg[07:00] <= tx_header_error_191_128_default[07:00];
      end
     else if (1'b1) begin
         tx_header_error_191_128_reg[07:00] <= i_tx_header_error_191_128_load_data[07:00];
       end
   end


// *****************************************************
// assign the register net to all the bits.
// *****************************************************
assign mmio_tx_header_error_191_128_wire = {
  tx_header_error_191_128_reg[63]    , tx_header_error_191_128_reg[62]    , tx_header_error_191_128_reg[61]    , tx_header_error_191_128_reg[60]    
, tx_header_error_191_128_reg[59]    , tx_header_error_191_128_reg[58]    , tx_header_error_191_128_reg[57]    , tx_header_error_191_128_reg[56]    
, tx_header_error_191_128_reg[55]    , tx_header_error_191_128_reg[54]    , tx_header_error_191_128_reg[53]    , tx_header_error_191_128_reg[52]    
, tx_header_error_191_128_reg[51]    , tx_header_error_191_128_reg[50]    , tx_header_error_191_128_reg[49]    , tx_header_error_191_128_reg[48]    
, tx_header_error_191_128_reg[47]    , tx_header_error_191_128_reg[46]    , tx_header_error_191_128_reg[45]    , tx_header_error_191_128_reg[44]    
, tx_header_error_191_128_reg[43]    , tx_header_error_191_128_reg[42]    , tx_header_error_191_128_reg[41]    , tx_header_error_191_128_reg[40]    
, tx_header_error_191_128_reg[39]    , tx_header_error_191_128_reg[38]    , tx_header_error_191_128_reg[37]    , tx_header_error_191_128_reg[36]    
, tx_header_error_191_128_reg[35]    , tx_header_error_191_128_reg[34]    , tx_header_error_191_128_reg[33]    , tx_header_error_191_128_reg[32]    
, tx_header_error_191_128_reg[31]    , tx_header_error_191_128_reg[30]    , tx_header_error_191_128_reg[29]    , tx_header_error_191_128_reg[28]    
, tx_header_error_191_128_reg[27]    , tx_header_error_191_128_reg[26]    , tx_header_error_191_128_reg[25]    , tx_header_error_191_128_reg[24]    
, tx_header_error_191_128_reg[23]    , tx_header_error_191_128_reg[22]    , tx_header_error_191_128_reg[21]    , tx_header_error_191_128_reg[20]    
, tx_header_error_191_128_reg[19]    , tx_header_error_191_128_reg[18]    , tx_header_error_191_128_reg[17]    , tx_header_error_191_128_reg[16]    
, tx_header_error_191_128_reg[15]    , tx_header_error_191_128_reg[14]    , tx_header_error_191_128_reg[13]    , tx_header_error_191_128_reg[12]    
, tx_header_error_191_128_reg[11]    , tx_header_error_191_128_reg[10]    , tx_header_error_191_128_reg[09]    , tx_header_error_191_128_reg[08]    
, tx_header_error_191_128_reg[07]    , tx_header_error_191_128_reg[06]    , tx_header_error_191_128_reg[05]    , tx_header_error_191_128_reg[04]    
, tx_header_error_191_128_reg[03]    , tx_header_error_191_128_reg[02]    , tx_header_error_191_128_reg[01]    , tx_header_error_191_128_reg[00]    };

// ******************************************************
// Register 0x048 mmio_tx_header_error_127_64
// ******************************************************
// ******************************************************
// Bit(s) 63:00 (tx_header_error_127_64) of Register 0x048 mmio_tx_header_error_127_64
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         tx_header_error_127_64_reg[63:56] <= tx_header_error_127_64_default[63:56];
      end
     else if (1'b1) begin
         tx_header_error_127_64_reg[63:56] <= i_tx_header_error_127_64_load_data[63:56];
       end
   end

// ******************************************************
// Bit(s) 63:00 (tx_header_error_127_64) of Register 0x048 mmio_tx_header_error_127_64
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         tx_header_error_127_64_reg[55:48] <= tx_header_error_127_64_default[55:48];
      end
     else if (1'b1) begin
         tx_header_error_127_64_reg[55:48] <= i_tx_header_error_127_64_load_data[55:48];
       end
   end

// ******************************************************
// Bit(s) 63:00 (tx_header_error_127_64) of Register 0x048 mmio_tx_header_error_127_64
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         tx_header_error_127_64_reg[47:40] <= tx_header_error_127_64_default[47:40];
      end
     else if (1'b1) begin
         tx_header_error_127_64_reg[47:40] <= i_tx_header_error_127_64_load_data[47:40];
       end
   end

// ******************************************************
// Bit(s) 63:00 (tx_header_error_127_64) of Register 0x048 mmio_tx_header_error_127_64
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         tx_header_error_127_64_reg[39:32] <= tx_header_error_127_64_default[39:32];
      end
     else if (1'b1) begin
         tx_header_error_127_64_reg[39:32] <= i_tx_header_error_127_64_load_data[39:32];
       end
   end

// ******************************************************
// Bit(s) 63:00 (tx_header_error_127_64) of Register 0x048 mmio_tx_header_error_127_64
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         tx_header_error_127_64_reg[31:24] <= tx_header_error_127_64_default[31:24];
      end
     else if (1'b1) begin
         tx_header_error_127_64_reg[31:24] <= i_tx_header_error_127_64_load_data[31:24];
       end
   end

// ******************************************************
// Bit(s) 63:00 (tx_header_error_127_64) of Register 0x048 mmio_tx_header_error_127_64
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         tx_header_error_127_64_reg[23:16] <= tx_header_error_127_64_default[23:16];
      end
     else if (1'b1) begin
         tx_header_error_127_64_reg[23:16] <= i_tx_header_error_127_64_load_data[23:16];
       end
   end

// ******************************************************
// Bit(s) 63:00 (tx_header_error_127_64) of Register 0x048 mmio_tx_header_error_127_64
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         tx_header_error_127_64_reg[15:08] <= tx_header_error_127_64_default[15:08];
      end
     else if (1'b1) begin
         tx_header_error_127_64_reg[15:08] <= i_tx_header_error_127_64_load_data[15:08];
       end
   end

// ******************************************************
// Bit(s) 63:00 (tx_header_error_127_64) of Register 0x048 mmio_tx_header_error_127_64
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         tx_header_error_127_64_reg[07:00] <= tx_header_error_127_64_default[07:00];
      end
     else if (1'b1) begin
         tx_header_error_127_64_reg[07:00] <= i_tx_header_error_127_64_load_data[07:00];
       end
   end


// *****************************************************
// assign the register net to all the bits.
// *****************************************************
assign mmio_tx_header_error_127_64_wire = {
  tx_header_error_127_64_reg[63]     , tx_header_error_127_64_reg[62]     , tx_header_error_127_64_reg[61]     , tx_header_error_127_64_reg[60]     
, tx_header_error_127_64_reg[59]     , tx_header_error_127_64_reg[58]     , tx_header_error_127_64_reg[57]     , tx_header_error_127_64_reg[56]     
, tx_header_error_127_64_reg[55]     , tx_header_error_127_64_reg[54]     , tx_header_error_127_64_reg[53]     , tx_header_error_127_64_reg[52]     
, tx_header_error_127_64_reg[51]     , tx_header_error_127_64_reg[50]     , tx_header_error_127_64_reg[49]     , tx_header_error_127_64_reg[48]     
, tx_header_error_127_64_reg[47]     , tx_header_error_127_64_reg[46]     , tx_header_error_127_64_reg[45]     , tx_header_error_127_64_reg[44]     
, tx_header_error_127_64_reg[43]     , tx_header_error_127_64_reg[42]     , tx_header_error_127_64_reg[41]     , tx_header_error_127_64_reg[40]     
, tx_header_error_127_64_reg[39]     , tx_header_error_127_64_reg[38]     , tx_header_error_127_64_reg[37]     , tx_header_error_127_64_reg[36]     
, tx_header_error_127_64_reg[35]     , tx_header_error_127_64_reg[34]     , tx_header_error_127_64_reg[33]     , tx_header_error_127_64_reg[32]     
, tx_header_error_127_64_reg[31]     , tx_header_error_127_64_reg[30]     , tx_header_error_127_64_reg[29]     , tx_header_error_127_64_reg[28]     
, tx_header_error_127_64_reg[27]     , tx_header_error_127_64_reg[26]     , tx_header_error_127_64_reg[25]     , tx_header_error_127_64_reg[24]     
, tx_header_error_127_64_reg[23]     , tx_header_error_127_64_reg[22]     , tx_header_error_127_64_reg[21]     , tx_header_error_127_64_reg[20]     
, tx_header_error_127_64_reg[19]     , tx_header_error_127_64_reg[18]     , tx_header_error_127_64_reg[17]     , tx_header_error_127_64_reg[16]     
, tx_header_error_127_64_reg[15]     , tx_header_error_127_64_reg[14]     , tx_header_error_127_64_reg[13]     , tx_header_error_127_64_reg[12]     
, tx_header_error_127_64_reg[11]     , tx_header_error_127_64_reg[10]     , tx_header_error_127_64_reg[09]     , tx_header_error_127_64_reg[08]     
, tx_header_error_127_64_reg[07]     , tx_header_error_127_64_reg[06]     , tx_header_error_127_64_reg[05]     , tx_header_error_127_64_reg[04]     
, tx_header_error_127_64_reg[03]     , tx_header_error_127_64_reg[02]     , tx_header_error_127_64_reg[01]     , tx_header_error_127_64_reg[00]     };

// ******************************************************
// Register 0x050 mmio_tx_header_error_63_00
// ******************************************************
// ******************************************************
// Bit(s) 63:00 (tx_header_error_63_00) of Register 0x050 mmio_tx_header_error_63_00
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         tx_header_error_63_00_reg[63:56] <= tx_header_error_63_00_default[63:56];
      end
     else if (1'b1) begin
         tx_header_error_63_00_reg[63:56] <= i_tx_header_error_63_00_load_data[63:56];
       end
   end

// ******************************************************
// Bit(s) 63:00 (tx_header_error_63_00) of Register 0x050 mmio_tx_header_error_63_00
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         tx_header_error_63_00_reg[55:48] <= tx_header_error_63_00_default[55:48];
      end
     else if (1'b1) begin
         tx_header_error_63_00_reg[55:48] <= i_tx_header_error_63_00_load_data[55:48];
       end
   end

// ******************************************************
// Bit(s) 63:00 (tx_header_error_63_00) of Register 0x050 mmio_tx_header_error_63_00
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         tx_header_error_63_00_reg[47:40] <= tx_header_error_63_00_default[47:40];
      end
     else if (1'b1) begin
         tx_header_error_63_00_reg[47:40] <= i_tx_header_error_63_00_load_data[47:40];
       end
   end

// ******************************************************
// Bit(s) 63:00 (tx_header_error_63_00) of Register 0x050 mmio_tx_header_error_63_00
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         tx_header_error_63_00_reg[39:32] <= tx_header_error_63_00_default[39:32];
      end
     else if (1'b1) begin
         tx_header_error_63_00_reg[39:32] <= i_tx_header_error_63_00_load_data[39:32];
       end
   end

// ******************************************************
// Bit(s) 63:00 (tx_header_error_63_00) of Register 0x050 mmio_tx_header_error_63_00
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         tx_header_error_63_00_reg[31:24] <= tx_header_error_63_00_default[31:24];
      end
     else if (1'b1) begin
         tx_header_error_63_00_reg[31:24] <= i_tx_header_error_63_00_load_data[31:24];
       end
   end

// ******************************************************
// Bit(s) 63:00 (tx_header_error_63_00) of Register 0x050 mmio_tx_header_error_63_00
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         tx_header_error_63_00_reg[23:16] <= tx_header_error_63_00_default[23:16];
      end
     else if (1'b1) begin
         tx_header_error_63_00_reg[23:16] <= i_tx_header_error_63_00_load_data[23:16];
       end
   end

// ******************************************************
// Bit(s) 63:00 (tx_header_error_63_00) of Register 0x050 mmio_tx_header_error_63_00
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         tx_header_error_63_00_reg[15:08] <= tx_header_error_63_00_default[15:08];
      end
     else if (1'b1) begin
         tx_header_error_63_00_reg[15:08] <= i_tx_header_error_63_00_load_data[15:08];
       end
   end

// ******************************************************
// Bit(s) 63:00 (tx_header_error_63_00) of Register 0x050 mmio_tx_header_error_63_00
// ******************************************************
   always @(posedge clk_csr) begin
      if (~pwr_good_csr_clk_n) begin
         tx_header_error_63_00_reg[07:00] <= tx_header_error_63_00_default[07:00];
      end
     else if (1'b1) begin
         tx_header_error_63_00_reg[07:00] <= i_tx_header_error_63_00_load_data[07:00];
       end
   end


// *****************************************************
// assign the register net to all the bits.
// *****************************************************
assign mmio_tx_header_error_63_00_wire = {
  tx_header_error_63_00_reg[63]      , tx_header_error_63_00_reg[62]      , tx_header_error_63_00_reg[61]      , tx_header_error_63_00_reg[60]      
, tx_header_error_63_00_reg[59]      , tx_header_error_63_00_reg[58]      , tx_header_error_63_00_reg[57]      , tx_header_error_63_00_reg[56]      
, tx_header_error_63_00_reg[55]      , tx_header_error_63_00_reg[54]      , tx_header_error_63_00_reg[53]      , tx_header_error_63_00_reg[52]      
, tx_header_error_63_00_reg[51]      , tx_header_error_63_00_reg[50]      , tx_header_error_63_00_reg[49]      , tx_header_error_63_00_reg[48]      
, tx_header_error_63_00_reg[47]      , tx_header_error_63_00_reg[46]      , tx_header_error_63_00_reg[45]      , tx_header_error_63_00_reg[44]      
, tx_header_error_63_00_reg[43]      , tx_header_error_63_00_reg[42]      , tx_header_error_63_00_reg[41]      , tx_header_error_63_00_reg[40]      
, tx_header_error_63_00_reg[39]      , tx_header_error_63_00_reg[38]      , tx_header_error_63_00_reg[37]      , tx_header_error_63_00_reg[36]      
, tx_header_error_63_00_reg[35]      , tx_header_error_63_00_reg[34]      , tx_header_error_63_00_reg[33]      , tx_header_error_63_00_reg[32]      
, tx_header_error_63_00_reg[31]      , tx_header_error_63_00_reg[30]      , tx_header_error_63_00_reg[29]      , tx_header_error_63_00_reg[28]      
, tx_header_error_63_00_reg[27]      , tx_header_error_63_00_reg[26]      , tx_header_error_63_00_reg[25]      , tx_header_error_63_00_reg[24]      
, tx_header_error_63_00_reg[23]      , tx_header_error_63_00_reg[22]      , tx_header_error_63_00_reg[21]      , tx_header_error_63_00_reg[20]      
, tx_header_error_63_00_reg[19]      , tx_header_error_63_00_reg[18]      , tx_header_error_63_00_reg[17]      , tx_header_error_63_00_reg[16]      
, tx_header_error_63_00_reg[15]      , tx_header_error_63_00_reg[14]      , tx_header_error_63_00_reg[13]      , tx_header_error_63_00_reg[12]      
, tx_header_error_63_00_reg[11]      , tx_header_error_63_00_reg[10]      , tx_header_error_63_00_reg[09]      , tx_header_error_63_00_reg[08]      
, tx_header_error_63_00_reg[07]      , tx_header_error_63_00_reg[06]      , tx_header_error_63_00_reg[05]      , tx_header_error_63_00_reg[04]      
, tx_header_error_63_00_reg[03]      , tx_header_error_63_00_reg[02]      , tx_header_error_63_00_reg[01]      , tx_header_error_63_00_reg[00]      };

// *****************************************************
// RTL for the first level muxes.
// *****************************************************
  always @(posedge clk_csr) begin
      csr_decode_mux_r4 <= 64'h00000000 // 0xff8
            | afu_intf_dfh_wire                   & {64{afu_intf_dfh_en_r3}}            // 0x000
            | afu_intf_scratchpad_wire            & {64{afu_intf_scratchpad_en_r3}}     // 0x008
            | afu_intf_error_wire                 & {64{afu_intf_error_en_r3}}          // 0x010
            | afu_intf_first_error_wire           & {64{afu_intf_first_error_en_r3}}    // 0x018
            | mmio_timeout_addr_wire              & {64{mmio_timeout_addr_en_r3}}       // 0x020
            | mmio_timeout_info_wire              & {64{mmio_timeout_info_en_r3}}       // 0x028
            | mmio_immediate_frozen_reg_wire      & {64{mmio_immediate_frozen_reg_en_r3}} // 0x030
            | mmio_tx_header_error_255_192_wire   & {64{mmio_tx_header_error_255_192_en_r3}} // 0x038
            | mmio_tx_header_error_191_128_wire   & {64{mmio_tx_header_error_191_128_en_r3}} // 0x040
            | mmio_tx_header_error_127_64_wire    & {64{mmio_tx_header_error_127_64_en_r3}} // 0x048
            | mmio_tx_header_error_63_00_wire     & {64{mmio_tx_header_error_63_00_en_r3}} // 0x050
              ;
    end

// *****************************************************
// Now onto everything on the clk clock domain.
// *****************************************************
   // *****************************************************
   // RTL for the final read mux (just an or gate) async signals masked by targeting_clkX_domain_register
   // *****************************************************
   always @(posedge clk_csr) begin
      csr_readdata <= csr_decode_mux_r4                                                          ; // 0xff8;
   end

   
   // synopsys translate_off
   //   wire [HI_ADDR_BIT:0] csr_address_real = {1'b1, csr_address, 2'h0};
   //`ifdef loggers_on
   //   
   //   always @(posedge clk_csr) begin
   //      if (csr_read & ~csr_waitrequest) begin
   //       $display("T:%8d INFO: %m RB RD addr:%x data:%x", $time, csr_address_real, csr_readdata);
   
   //      end
   //      if (csr_write & ~csr_waitrequest) begin
   //       $display("T:%8d INFO: %m RB WR addr:%x data:%x", $time, csr_address_real, csr_wdata);
   //      end
   //   end
   //`endif
   // synopsys translate_on
   
endmodule
