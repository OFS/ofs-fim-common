// Copyright (C) 2023 Intel Corporation
// SPDX-License-Identifier: MIT

/**
 * Abstract:
 * Defines a virtual sequencer for the testbench ENV.  This sequencer obtains
 * a handle to the reset interface using the config db.  This allows
 * reset sequences to be written for this sequencer.
 */

`ifndef GUARD_pf_vf_mux_virtual_sequencer_SV
`define GUARD_pf_vf_mux_virtual_sequencer_SV

class pf_vf_mux_virtual_sequencer extends uvm_sequencer;

  /** Typedef of the reset modport to simplify access */
  typedef virtual axi_reset_if.axi_reset_modport AXI_RESET_MP;

  /** Reset modport provides access to the reset signal */
  AXI_RESET_MP reset_mp;

  `uvm_component_utils(pf_vf_mux_virtual_sequencer)
   svt_axi_master_sequencer    master_sequencer_H;
   svt_axi_master_sequencer    master_sequencer_D0;
   svt_axi_master_sequencer    master_sequencer_D1;
   svt_axi_master_sequencer    master_sequencer_D2;
   svt_axi_master_sequencer    master_sequencer_D3;
   svt_axi_master_sequencer    master_sequencer_D4;
   svt_axi_master_sequencer    master_sequencer_D5;
   svt_axi_master_sequencer    master_sequencer_D6;
   svt_axi_master_sequencer    master_sequencer_D7;
   svt_axi_master_sequencer    master_sequencer_D8;
   svt_axi_master_sequencer    master_sequencer_D9;
   svt_axi_master_sequencer    master_sequencer_D10;
   svt_axi_master_sequencer    master_sequencer_D11;
   svt_axi_master_sequencer    master_sequencer_D12;
   svt_axi_master_sequencer    master_sequencer_D13;
   svt_axi_master_sequencer    master_sequencer_D14;
   svt_axi_master_sequencer    master_sequencer_D15;
   svt_axi_master_sequencer    master_sequencer_DN0;
   svt_axi_master_sequencer    master_sequencer_DN1;
   svt_axi_master_sequencer    master_sequencer_DN2;
   svt_axi_master_sequencer    master_sequencer_DN3;
   svt_axi_master_sequencer    master_sequencer_DN4;
   svt_axi_master_sequencer    master_sequencer_DN5;
   svt_axi_master_sequencer    master_sequencer_DN6;
   svt_axi_master_sequencer    master_sequencer_DN7;
   svt_axi_master_sequencer    master_sequencer_DN8;
   svt_axi_master_sequencer    master_sequencer_DN9;
   svt_axi_master_sequencer    master_sequencer_DN10;
   svt_axi_master_sequencer    master_sequencer_DN11;
   svt_axi_master_sequencer    master_sequencer_DN12;
   svt_axi_master_sequencer    master_sequencer_DN13;
   svt_axi_master_sequencer    master_sequencer_DN14;
   svt_axi_master_sequencer    master_sequencer_DN15;
   `ifdef TB_CONFIG_4
   svt_axi_master_sequencer    master_sequencer_D16;
   svt_axi_master_sequencer    master_sequencer_D17;
   svt_axi_master_sequencer    master_sequencer_D18;
   svt_axi_master_sequencer    master_sequencer_D19;
   svt_axi_master_sequencer    master_sequencer_D20;
   svt_axi_master_sequencer    master_sequencer_D21;
   svt_axi_master_sequencer    master_sequencer_D22;
   svt_axi_master_sequencer    master_sequencer_D23;
   svt_axi_master_sequencer    master_sequencer_D24;
   svt_axi_master_sequencer    master_sequencer_D25;
   svt_axi_master_sequencer    master_sequencer_D26;
   svt_axi_master_sequencer    master_sequencer_D27;
   svt_axi_master_sequencer    master_sequencer_D28;
   svt_axi_master_sequencer    master_sequencer_D29;
   svt_axi_master_sequencer    master_sequencer_D30;
   svt_axi_master_sequencer    master_sequencer_D31;
   svt_axi_master_sequencer    master_sequencer_D32;
   svt_axi_master_sequencer    master_sequencer_D33;
   svt_axi_master_sequencer    master_sequencer_D34;
   svt_axi_master_sequencer    master_sequencer_D35;
   svt_axi_master_sequencer    master_sequencer_D36;
   svt_axi_master_sequencer    master_sequencer_D37;
   svt_axi_master_sequencer    master_sequencer_D38;
   svt_axi_master_sequencer    master_sequencer_D39;
   svt_axi_master_sequencer    master_sequencer_D40;
   svt_axi_master_sequencer    master_sequencer_D41;
   svt_axi_master_sequencer    master_sequencer_D42;
   svt_axi_master_sequencer    master_sequencer_D43;
   svt_axi_master_sequencer    master_sequencer_D44;
   svt_axi_master_sequencer    master_sequencer_D45;
   svt_axi_master_sequencer    master_sequencer_D46;
   svt_axi_master_sequencer    master_sequencer_D47;
   svt_axi_master_sequencer    master_sequencer_D48;
   svt_axi_master_sequencer    master_sequencer_D49;
   svt_axi_master_sequencer    master_sequencer_D50;
   svt_axi_master_sequencer    master_sequencer_D51;
   svt_axi_master_sequencer    master_sequencer_D52;
   svt_axi_master_sequencer    master_sequencer_D53;
   svt_axi_master_sequencer    master_sequencer_D54;
   svt_axi_master_sequencer    master_sequencer_D55;
   svt_axi_master_sequencer    master_sequencer_D56;
   svt_axi_master_sequencer    master_sequencer_D57;
   svt_axi_master_sequencer    master_sequencer_D58;
   svt_axi_master_sequencer    master_sequencer_D59;
   svt_axi_master_sequencer    master_sequencer_D60;
   svt_axi_master_sequencer    master_sequencer_D61;
   svt_axi_master_sequencer    master_sequencer_D62;
   svt_axi_master_sequencer    master_sequencer_D63;
   svt_axi_master_sequencer    master_sequencer_D64;
   svt_axi_master_sequencer    master_sequencer_D65;
   svt_axi_master_sequencer    master_sequencer_D66;
   svt_axi_master_sequencer    master_sequencer_D67;
   svt_axi_master_sequencer    master_sequencer_D68;
   svt_axi_master_sequencer    master_sequencer_D69;
   svt_axi_master_sequencer    master_sequencer_D70;
   svt_axi_master_sequencer    master_sequencer_D71;
   svt_axi_master_sequencer    master_sequencer_D72;
   svt_axi_master_sequencer    master_sequencer_D73;
   svt_axi_master_sequencer    master_sequencer_D74;
   svt_axi_master_sequencer    master_sequencer_D75;
   svt_axi_master_sequencer    master_sequencer_D76;
   svt_axi_master_sequencer    master_sequencer_D77;
   svt_axi_master_sequencer    master_sequencer_D78;
   svt_axi_master_sequencer    master_sequencer_D79;
   svt_axi_master_sequencer    master_sequencer_D80;
   svt_axi_master_sequencer    master_sequencer_D81;
   svt_axi_master_sequencer    master_sequencer_D82;
   svt_axi_master_sequencer    master_sequencer_D83;
   svt_axi_master_sequencer    master_sequencer_D84;
   svt_axi_master_sequencer    master_sequencer_D85;
   svt_axi_master_sequencer    master_sequencer_D86;
   svt_axi_master_sequencer    master_sequencer_D87;
   svt_axi_master_sequencer    master_sequencer_D88;
   svt_axi_master_sequencer    master_sequencer_D89;
   svt_axi_master_sequencer    master_sequencer_D90;
   svt_axi_master_sequencer    master_sequencer_D91;
   svt_axi_master_sequencer    master_sequencer_D92;
   svt_axi_master_sequencer    master_sequencer_D93;
   svt_axi_master_sequencer    master_sequencer_D94;
   svt_axi_master_sequencer    master_sequencer_D95;
   svt_axi_master_sequencer    master_sequencer_D96;
   svt_axi_master_sequencer    master_sequencer_D97;
   svt_axi_master_sequencer    master_sequencer_D98;
   svt_axi_master_sequencer    master_sequencer_D99;
   svt_axi_master_sequencer    master_sequencer_D100;
   svt_axi_master_sequencer    master_sequencer_D101;
   svt_axi_master_sequencer    master_sequencer_D102;
   svt_axi_master_sequencer    master_sequencer_D103;
   svt_axi_master_sequencer    master_sequencer_D104;
   svt_axi_master_sequencer    master_sequencer_D105;
   svt_axi_master_sequencer    master_sequencer_D106;
   svt_axi_master_sequencer    master_sequencer_D107;
   svt_axi_master_sequencer    master_sequencer_D108;
   svt_axi_master_sequencer    master_sequencer_D109;
   svt_axi_master_sequencer    master_sequencer_D110;
   svt_axi_master_sequencer    master_sequencer_D111;
   svt_axi_master_sequencer    master_sequencer_D112;
   svt_axi_master_sequencer    master_sequencer_D113;
   svt_axi_master_sequencer    master_sequencer_D114;
   svt_axi_master_sequencer    master_sequencer_D115;
   svt_axi_master_sequencer    master_sequencer_D116;
   svt_axi_master_sequencer    master_sequencer_D117;
   svt_axi_master_sequencer    master_sequencer_D118;
   svt_axi_master_sequencer    master_sequencer_D119;
   svt_axi_master_sequencer    master_sequencer_D120;
   svt_axi_master_sequencer    master_sequencer_D121;
   svt_axi_master_sequencer    master_sequencer_D122;
   svt_axi_master_sequencer    master_sequencer_D123;
   svt_axi_master_sequencer    master_sequencer_D124;
   svt_axi_master_sequencer    master_sequencer_D125;
   svt_axi_master_sequencer    master_sequencer_D126;
   svt_axi_master_sequencer    master_sequencer_D127;
   svt_axi_master_sequencer    master_sequencer_D128;
   svt_axi_master_sequencer    master_sequencer_D129;
   svt_axi_master_sequencer    master_sequencer_D130;
   svt_axi_master_sequencer    master_sequencer_D131;
   svt_axi_master_sequencer    master_sequencer_D132;
   svt_axi_master_sequencer    master_sequencer_D133;
   svt_axi_master_sequencer    master_sequencer_D134;
   svt_axi_master_sequencer    master_sequencer_D135;
   svt_axi_master_sequencer    master_sequencer_D136;
   svt_axi_master_sequencer    master_sequencer_D137;
   svt_axi_master_sequencer    master_sequencer_D138;
   svt_axi_master_sequencer    master_sequencer_D139;
   svt_axi_master_sequencer    master_sequencer_D140;
   svt_axi_master_sequencer    master_sequencer_D141;
   svt_axi_master_sequencer    master_sequencer_D142;
   svt_axi_master_sequencer    master_sequencer_D143;
   svt_axi_master_sequencer    master_sequencer_D144;
   svt_axi_master_sequencer    master_sequencer_D145;
   svt_axi_master_sequencer    master_sequencer_D146;
   svt_axi_master_sequencer    master_sequencer_D147;
   svt_axi_master_sequencer    master_sequencer_D148;
   svt_axi_master_sequencer    master_sequencer_D149;
   svt_axi_master_sequencer    master_sequencer_D150;
   svt_axi_master_sequencer    master_sequencer_D151;
   svt_axi_master_sequencer    master_sequencer_D152;
   svt_axi_master_sequencer    master_sequencer_D153;
   svt_axi_master_sequencer    master_sequencer_D154;
   svt_axi_master_sequencer    master_sequencer_D155;
   svt_axi_master_sequencer    master_sequencer_D156;
   svt_axi_master_sequencer    master_sequencer_D157;
   svt_axi_master_sequencer    master_sequencer_D158;
   svt_axi_master_sequencer    master_sequencer_D159;
   svt_axi_master_sequencer    master_sequencer_D160;
   svt_axi_master_sequencer    master_sequencer_D161;
   svt_axi_master_sequencer    master_sequencer_D162;
   svt_axi_master_sequencer    master_sequencer_D163;
   svt_axi_master_sequencer    master_sequencer_D164;
   svt_axi_master_sequencer    master_sequencer_D165;
   svt_axi_master_sequencer    master_sequencer_D166;
   svt_axi_master_sequencer    master_sequencer_D167;
   svt_axi_master_sequencer    master_sequencer_D168;
   svt_axi_master_sequencer    master_sequencer_D169;
   svt_axi_master_sequencer    master_sequencer_D170;
   svt_axi_master_sequencer    master_sequencer_D171;
   svt_axi_master_sequencer    master_sequencer_D172;
   svt_axi_master_sequencer    master_sequencer_D173;
   svt_axi_master_sequencer    master_sequencer_D174;
   svt_axi_master_sequencer    master_sequencer_D175;
   svt_axi_master_sequencer    master_sequencer_D176;
   svt_axi_master_sequencer    master_sequencer_D177;
   svt_axi_master_sequencer    master_sequencer_D178;
   svt_axi_master_sequencer    master_sequencer_D179;
   svt_axi_master_sequencer    master_sequencer_D180;
   svt_axi_master_sequencer    master_sequencer_D181;
   svt_axi_master_sequencer    master_sequencer_D182;
   svt_axi_master_sequencer    master_sequencer_D183;
   svt_axi_master_sequencer    master_sequencer_D184;
   svt_axi_master_sequencer    master_sequencer_D185;
   svt_axi_master_sequencer    master_sequencer_D186;
   svt_axi_master_sequencer    master_sequencer_D187;
   svt_axi_master_sequencer    master_sequencer_D188;
   svt_axi_master_sequencer    master_sequencer_D189;
   svt_axi_master_sequencer    master_sequencer_D190;
   svt_axi_master_sequencer    master_sequencer_D191;
   svt_axi_master_sequencer    master_sequencer_D192;
   svt_axi_master_sequencer    master_sequencer_D193;
   svt_axi_master_sequencer    master_sequencer_D194;
   svt_axi_master_sequencer    master_sequencer_D195;
   svt_axi_master_sequencer    master_sequencer_D196;
   svt_axi_master_sequencer    master_sequencer_D197;
   svt_axi_master_sequencer    master_sequencer_D198;
   svt_axi_master_sequencer    master_sequencer_D199;
   svt_axi_master_sequencer    master_sequencer_D200;
   svt_axi_master_sequencer    master_sequencer_D201;
   svt_axi_master_sequencer    master_sequencer_D202;
   svt_axi_master_sequencer    master_sequencer_D203;
   svt_axi_master_sequencer    master_sequencer_D204;
   svt_axi_master_sequencer    master_sequencer_D205;
   svt_axi_master_sequencer    master_sequencer_D206;
   svt_axi_master_sequencer    master_sequencer_D207;
   svt_axi_master_sequencer    master_sequencer_D208;
   svt_axi_master_sequencer    master_sequencer_D209;
   svt_axi_master_sequencer    master_sequencer_D210;
   svt_axi_master_sequencer    master_sequencer_D211;
   svt_axi_master_sequencer    master_sequencer_D212;
   svt_axi_master_sequencer    master_sequencer_D213;
   svt_axi_master_sequencer    master_sequencer_D214;
   svt_axi_master_sequencer    master_sequencer_D215;
   svt_axi_master_sequencer    master_sequencer_D216;
   svt_axi_master_sequencer    master_sequencer_D217;
   svt_axi_master_sequencer    master_sequencer_D218;
   svt_axi_master_sequencer    master_sequencer_D219;
   svt_axi_master_sequencer    master_sequencer_D220;
   svt_axi_master_sequencer    master_sequencer_D221;
   svt_axi_master_sequencer    master_sequencer_D222;
   svt_axi_master_sequencer    master_sequencer_D223;
   svt_axi_master_sequencer    master_sequencer_D224;
   svt_axi_master_sequencer    master_sequencer_D225;
   svt_axi_master_sequencer    master_sequencer_D226;
   svt_axi_master_sequencer    master_sequencer_D227;
   svt_axi_master_sequencer    master_sequencer_D228;
   svt_axi_master_sequencer    master_sequencer_D229;
   svt_axi_master_sequencer    master_sequencer_D230;
   svt_axi_master_sequencer    master_sequencer_D231;
   svt_axi_master_sequencer    master_sequencer_D232;
   svt_axi_master_sequencer    master_sequencer_D233;
   svt_axi_master_sequencer    master_sequencer_D234;
   svt_axi_master_sequencer    master_sequencer_D235;
   svt_axi_master_sequencer    master_sequencer_D236;
   svt_axi_master_sequencer    master_sequencer_D237;
   svt_axi_master_sequencer    master_sequencer_D238;
   svt_axi_master_sequencer    master_sequencer_D239;
   svt_axi_master_sequencer    master_sequencer_D240;
   svt_axi_master_sequencer    master_sequencer_D241;
   svt_axi_master_sequencer    master_sequencer_D242;
   svt_axi_master_sequencer    master_sequencer_D243;
   svt_axi_master_sequencer    master_sequencer_D244;
   svt_axi_master_sequencer    master_sequencer_D245;
   svt_axi_master_sequencer    master_sequencer_D246;
   svt_axi_master_sequencer    master_sequencer_D247;
   svt_axi_master_sequencer    master_sequencer_D248;
   svt_axi_master_sequencer    master_sequencer_D249;
   svt_axi_master_sequencer    master_sequencer_D250;
   svt_axi_master_sequencer    master_sequencer_D251;
   svt_axi_master_sequencer    master_sequencer_D252;
   svt_axi_master_sequencer    master_sequencer_D253;
   svt_axi_master_sequencer    master_sequencer_D254;
   svt_axi_master_sequencer    master_sequencer_D255;
   svt_axi_master_sequencer    master_sequencer_D256;
   svt_axi_master_sequencer    master_sequencer_D257;
   svt_axi_master_sequencer    master_sequencer_D258;
   svt_axi_master_sequencer    master_sequencer_D259;
   svt_axi_master_sequencer    master_sequencer_D260;
   svt_axi_master_sequencer    master_sequencer_D261;
   svt_axi_master_sequencer    master_sequencer_D262;
   svt_axi_master_sequencer    master_sequencer_D263;
   svt_axi_master_sequencer    master_sequencer_D264;
   svt_axi_master_sequencer    master_sequencer_D265;
   svt_axi_master_sequencer    master_sequencer_D266;
   svt_axi_master_sequencer    master_sequencer_D267;
   svt_axi_master_sequencer    master_sequencer_D268;
   svt_axi_master_sequencer    master_sequencer_D269;
   svt_axi_master_sequencer    master_sequencer_D270;
   svt_axi_master_sequencer    master_sequencer_D271;
   svt_axi_master_sequencer    master_sequencer_D272;
   svt_axi_master_sequencer    master_sequencer_D273;
   svt_axi_master_sequencer    master_sequencer_D274;
   svt_axi_master_sequencer    master_sequencer_D275;
   svt_axi_master_sequencer    master_sequencer_D276;
   svt_axi_master_sequencer    master_sequencer_D277;
   svt_axi_master_sequencer    master_sequencer_D278;
   svt_axi_master_sequencer    master_sequencer_D279;
   svt_axi_master_sequencer    master_sequencer_D280;
   svt_axi_master_sequencer    master_sequencer_D281;
   svt_axi_master_sequencer    master_sequencer_D282;
   svt_axi_master_sequencer    master_sequencer_D283;
   svt_axi_master_sequencer    master_sequencer_D284;
   svt_axi_master_sequencer    master_sequencer_D285;
   svt_axi_master_sequencer    master_sequencer_D286;
   svt_axi_master_sequencer    master_sequencer_D287;
   svt_axi_master_sequencer    master_sequencer_D288;
   svt_axi_master_sequencer    master_sequencer_D289;
   svt_axi_master_sequencer    master_sequencer_D290;
   svt_axi_master_sequencer    master_sequencer_D291;
   svt_axi_master_sequencer    master_sequencer_D292;
   svt_axi_master_sequencer    master_sequencer_D293;
   svt_axi_master_sequencer    master_sequencer_D294;
   svt_axi_master_sequencer    master_sequencer_D295;
   svt_axi_master_sequencer    master_sequencer_D296;
   svt_axi_master_sequencer    master_sequencer_D297;
   svt_axi_master_sequencer    master_sequencer_D298;
   svt_axi_master_sequencer    master_sequencer_D299;
   svt_axi_master_sequencer    master_sequencer_D300;
   svt_axi_master_sequencer    master_sequencer_D301;
   svt_axi_master_sequencer    master_sequencer_D302;
   svt_axi_master_sequencer    master_sequencer_D303;
   svt_axi_master_sequencer    master_sequencer_D304;
   svt_axi_master_sequencer    master_sequencer_D305;
   svt_axi_master_sequencer    master_sequencer_D306;
   svt_axi_master_sequencer    master_sequencer_D307;
   svt_axi_master_sequencer    master_sequencer_D308;
   svt_axi_master_sequencer    master_sequencer_D309;
   svt_axi_master_sequencer    master_sequencer_D310;
   svt_axi_master_sequencer    master_sequencer_D311;
   svt_axi_master_sequencer    master_sequencer_D312;
   svt_axi_master_sequencer    master_sequencer_D313;
   svt_axi_master_sequencer    master_sequencer_D314;
   svt_axi_master_sequencer    master_sequencer_D315;
   svt_axi_master_sequencer    master_sequencer_D316;
   svt_axi_master_sequencer    master_sequencer_D317;
   svt_axi_master_sequencer    master_sequencer_D318;
   svt_axi_master_sequencer    master_sequencer_D319;
   svt_axi_master_sequencer    master_sequencer_D320;
   svt_axi_master_sequencer    master_sequencer_D321;
   svt_axi_master_sequencer    master_sequencer_D322;
   svt_axi_master_sequencer    master_sequencer_D323;
   svt_axi_master_sequencer    master_sequencer_D324;
   svt_axi_master_sequencer    master_sequencer_D325;
   svt_axi_master_sequencer    master_sequencer_D326;
   svt_axi_master_sequencer    master_sequencer_D327;
   svt_axi_master_sequencer    master_sequencer_D328;
   svt_axi_master_sequencer    master_sequencer_D329;
   svt_axi_master_sequencer    master_sequencer_D330;
   svt_axi_master_sequencer    master_sequencer_D331;
   svt_axi_master_sequencer    master_sequencer_D332;
   svt_axi_master_sequencer    master_sequencer_D333;
   svt_axi_master_sequencer    master_sequencer_D334;
   svt_axi_master_sequencer    master_sequencer_D335;
   svt_axi_master_sequencer    master_sequencer_D336;
   svt_axi_master_sequencer    master_sequencer_D337;
   svt_axi_master_sequencer    master_sequencer_D338;
   svt_axi_master_sequencer    master_sequencer_D339;
   svt_axi_master_sequencer    master_sequencer_D340;
   svt_axi_master_sequencer    master_sequencer_D341;
   svt_axi_master_sequencer    master_sequencer_D342;
   svt_axi_master_sequencer    master_sequencer_D343;
   svt_axi_master_sequencer    master_sequencer_D344;
   svt_axi_master_sequencer    master_sequencer_D345;
   svt_axi_master_sequencer    master_sequencer_D346;
   svt_axi_master_sequencer    master_sequencer_D347;
   svt_axi_master_sequencer    master_sequencer_D348;
   svt_axi_master_sequencer    master_sequencer_D349;
   svt_axi_master_sequencer    master_sequencer_D350;
   svt_axi_master_sequencer    master_sequencer_D351;
   svt_axi_master_sequencer    master_sequencer_D352;
   svt_axi_master_sequencer    master_sequencer_D353;
   svt_axi_master_sequencer    master_sequencer_D354;
   svt_axi_master_sequencer    master_sequencer_D355;
   svt_axi_master_sequencer    master_sequencer_D356;
   svt_axi_master_sequencer    master_sequencer_D357;
   svt_axi_master_sequencer    master_sequencer_D358;
   svt_axi_master_sequencer    master_sequencer_D359;
   svt_axi_master_sequencer    master_sequencer_D360;
   svt_axi_master_sequencer    master_sequencer_D361;
   svt_axi_master_sequencer    master_sequencer_D362;
   svt_axi_master_sequencer    master_sequencer_D363;
   svt_axi_master_sequencer    master_sequencer_D364;
   svt_axi_master_sequencer    master_sequencer_D365;
   svt_axi_master_sequencer    master_sequencer_D366;
   svt_axi_master_sequencer    master_sequencer_D367;
   svt_axi_master_sequencer    master_sequencer_D368;
   svt_axi_master_sequencer    master_sequencer_D369;
   svt_axi_master_sequencer    master_sequencer_D370;
   svt_axi_master_sequencer    master_sequencer_D371;
   svt_axi_master_sequencer    master_sequencer_D372;
   svt_axi_master_sequencer    master_sequencer_D373;
   svt_axi_master_sequencer    master_sequencer_D374;
   svt_axi_master_sequencer    master_sequencer_D375;
   svt_axi_master_sequencer    master_sequencer_D376;
   svt_axi_master_sequencer    master_sequencer_D377;
   svt_axi_master_sequencer    master_sequencer_D378;
   svt_axi_master_sequencer    master_sequencer_D379;
   svt_axi_master_sequencer    master_sequencer_D380;
   svt_axi_master_sequencer    master_sequencer_D381;
   svt_axi_master_sequencer    master_sequencer_D382;
   svt_axi_master_sequencer    master_sequencer_D383;
   svt_axi_master_sequencer    master_sequencer_D384;
   svt_axi_master_sequencer    master_sequencer_D385;
   svt_axi_master_sequencer    master_sequencer_D386;
   svt_axi_master_sequencer    master_sequencer_D387;
   svt_axi_master_sequencer    master_sequencer_D388;
   svt_axi_master_sequencer    master_sequencer_D389;
   svt_axi_master_sequencer    master_sequencer_D390;
   svt_axi_master_sequencer    master_sequencer_D391;
   svt_axi_master_sequencer    master_sequencer_D392;
   svt_axi_master_sequencer    master_sequencer_D393;
   svt_axi_master_sequencer    master_sequencer_D394;
   svt_axi_master_sequencer    master_sequencer_D395;
   svt_axi_master_sequencer    master_sequencer_D396;
   svt_axi_master_sequencer    master_sequencer_D397;
   svt_axi_master_sequencer    master_sequencer_D398;
   svt_axi_master_sequencer    master_sequencer_D399;
   svt_axi_master_sequencer    master_sequencer_D400;
   svt_axi_master_sequencer    master_sequencer_D401;
   svt_axi_master_sequencer    master_sequencer_D402;
   svt_axi_master_sequencer    master_sequencer_D403;
   svt_axi_master_sequencer    master_sequencer_D404;
   svt_axi_master_sequencer    master_sequencer_D405;
   svt_axi_master_sequencer    master_sequencer_D406;
   svt_axi_master_sequencer    master_sequencer_D407;
   svt_axi_master_sequencer    master_sequencer_D408;
   svt_axi_master_sequencer    master_sequencer_D409;
   svt_axi_master_sequencer    master_sequencer_D410;
   svt_axi_master_sequencer    master_sequencer_D411;
   svt_axi_master_sequencer    master_sequencer_D412;
   svt_axi_master_sequencer    master_sequencer_D413;
   svt_axi_master_sequencer    master_sequencer_D414;
   svt_axi_master_sequencer    master_sequencer_D415;
   svt_axi_master_sequencer    master_sequencer_D416;
   svt_axi_master_sequencer    master_sequencer_D417;
   svt_axi_master_sequencer    master_sequencer_D418;
   svt_axi_master_sequencer    master_sequencer_D419;
   svt_axi_master_sequencer    master_sequencer_D420;
   svt_axi_master_sequencer    master_sequencer_D421;
   svt_axi_master_sequencer    master_sequencer_D422;
   svt_axi_master_sequencer    master_sequencer_D423;
   svt_axi_master_sequencer    master_sequencer_D424;
   svt_axi_master_sequencer    master_sequencer_D425;
   svt_axi_master_sequencer    master_sequencer_D426;
   svt_axi_master_sequencer    master_sequencer_D427;
   svt_axi_master_sequencer    master_sequencer_D428;
   svt_axi_master_sequencer    master_sequencer_D429;
   svt_axi_master_sequencer    master_sequencer_D430;
   svt_axi_master_sequencer    master_sequencer_D431;
   svt_axi_master_sequencer    master_sequencer_D432;
   svt_axi_master_sequencer    master_sequencer_D433;
   svt_axi_master_sequencer    master_sequencer_D434;
   svt_axi_master_sequencer    master_sequencer_D435;
   svt_axi_master_sequencer    master_sequencer_D436;
   svt_axi_master_sequencer    master_sequencer_D437;
   svt_axi_master_sequencer    master_sequencer_D438;
   svt_axi_master_sequencer    master_sequencer_D439;
   svt_axi_master_sequencer    master_sequencer_D440;
   svt_axi_master_sequencer    master_sequencer_D441;
   svt_axi_master_sequencer    master_sequencer_D442;
   svt_axi_master_sequencer    master_sequencer_D443;
   svt_axi_master_sequencer    master_sequencer_D444;
   svt_axi_master_sequencer    master_sequencer_D445;
   svt_axi_master_sequencer    master_sequencer_D446;
   svt_axi_master_sequencer    master_sequencer_D447;
   svt_axi_master_sequencer    master_sequencer_D448;
   svt_axi_master_sequencer    master_sequencer_D449;
   svt_axi_master_sequencer    master_sequencer_D450;
   svt_axi_master_sequencer    master_sequencer_D451;
   svt_axi_master_sequencer    master_sequencer_D452;
   svt_axi_master_sequencer    master_sequencer_D453;
   svt_axi_master_sequencer    master_sequencer_D454;
   svt_axi_master_sequencer    master_sequencer_D455;
   svt_axi_master_sequencer    master_sequencer_D456;
   svt_axi_master_sequencer    master_sequencer_D457;
   svt_axi_master_sequencer    master_sequencer_D458;
   svt_axi_master_sequencer    master_sequencer_D459;
   svt_axi_master_sequencer    master_sequencer_D460;
   svt_axi_master_sequencer    master_sequencer_D461;
   svt_axi_master_sequencer    master_sequencer_D462;
   svt_axi_master_sequencer    master_sequencer_D463;
   svt_axi_master_sequencer    master_sequencer_D464;
   svt_axi_master_sequencer    master_sequencer_D465;
   svt_axi_master_sequencer    master_sequencer_D466;
   svt_axi_master_sequencer    master_sequencer_D467;
   svt_axi_master_sequencer    master_sequencer_D468;
   svt_axi_master_sequencer    master_sequencer_D469;
   svt_axi_master_sequencer    master_sequencer_D470;
   svt_axi_master_sequencer    master_sequencer_D471;
   svt_axi_master_sequencer    master_sequencer_D472;
   svt_axi_master_sequencer    master_sequencer_D473;
   svt_axi_master_sequencer    master_sequencer_D474;
   svt_axi_master_sequencer    master_sequencer_D475;
   svt_axi_master_sequencer    master_sequencer_D476;
   svt_axi_master_sequencer    master_sequencer_D477;
   svt_axi_master_sequencer    master_sequencer_D478;
   svt_axi_master_sequencer    master_sequencer_D479;
   svt_axi_master_sequencer    master_sequencer_D480;
   svt_axi_master_sequencer    master_sequencer_D481;
   svt_axi_master_sequencer    master_sequencer_D482;
   svt_axi_master_sequencer    master_sequencer_D483;
   svt_axi_master_sequencer    master_sequencer_D484;
   svt_axi_master_sequencer    master_sequencer_D485;
   svt_axi_master_sequencer    master_sequencer_D486;
   svt_axi_master_sequencer    master_sequencer_D487;
   svt_axi_master_sequencer    master_sequencer_D488;
   svt_axi_master_sequencer    master_sequencer_D489;
   svt_axi_master_sequencer    master_sequencer_D490;
   svt_axi_master_sequencer    master_sequencer_D491;
   svt_axi_master_sequencer    master_sequencer_D492;
   svt_axi_master_sequencer    master_sequencer_D493;
   svt_axi_master_sequencer    master_sequencer_D494;
   svt_axi_master_sequencer    master_sequencer_D495;
   svt_axi_master_sequencer    master_sequencer_D496;
   svt_axi_master_sequencer    master_sequencer_D497;
   svt_axi_master_sequencer    master_sequencer_D498;
   svt_axi_master_sequencer    master_sequencer_D499;
   svt_axi_master_sequencer    master_sequencer_D500;
   svt_axi_master_sequencer    master_sequencer_D501;
   svt_axi_master_sequencer    master_sequencer_D502;
   svt_axi_master_sequencer    master_sequencer_D503;
   svt_axi_master_sequencer    master_sequencer_D504;
   svt_axi_master_sequencer    master_sequencer_D505;
   svt_axi_master_sequencer    master_sequencer_D506;
   svt_axi_master_sequencer    master_sequencer_D507;
   svt_axi_master_sequencer    master_sequencer_D508;
   svt_axi_master_sequencer    master_sequencer_D509;
   svt_axi_master_sequencer    master_sequencer_D510;
   svt_axi_master_sequencer    master_sequencer_D511;
   svt_axi_master_sequencer    master_sequencer_D512;
   svt_axi_master_sequencer    master_sequencer_D513;
   svt_axi_master_sequencer    master_sequencer_D514;
   svt_axi_master_sequencer    master_sequencer_D515;
   svt_axi_master_sequencer    master_sequencer_D516;
   svt_axi_master_sequencer    master_sequencer_D517;
   svt_axi_master_sequencer    master_sequencer_D518;
   svt_axi_master_sequencer    master_sequencer_D519;
   svt_axi_master_sequencer    master_sequencer_D520;
   svt_axi_master_sequencer    master_sequencer_D521;
   svt_axi_master_sequencer    master_sequencer_D522;
   svt_axi_master_sequencer    master_sequencer_D523;
   svt_axi_master_sequencer    master_sequencer_D524;
   svt_axi_master_sequencer    master_sequencer_D525;
   svt_axi_master_sequencer    master_sequencer_D526;
   svt_axi_master_sequencer    master_sequencer_D527;
   svt_axi_master_sequencer    master_sequencer_D528;
   svt_axi_master_sequencer    master_sequencer_D529;
   svt_axi_master_sequencer    master_sequencer_D530;
   svt_axi_master_sequencer    master_sequencer_D531;
   svt_axi_master_sequencer    master_sequencer_D532;
   svt_axi_master_sequencer    master_sequencer_D533;
   svt_axi_master_sequencer    master_sequencer_D534;
   svt_axi_master_sequencer    master_sequencer_D535;
   svt_axi_master_sequencer    master_sequencer_D536;
   svt_axi_master_sequencer    master_sequencer_D537;
   svt_axi_master_sequencer    master_sequencer_D538;
   svt_axi_master_sequencer    master_sequencer_D539;
   svt_axi_master_sequencer    master_sequencer_D540;
   svt_axi_master_sequencer    master_sequencer_D541;
   svt_axi_master_sequencer    master_sequencer_D542;
   svt_axi_master_sequencer    master_sequencer_D543;
   svt_axi_master_sequencer    master_sequencer_D544;
   svt_axi_master_sequencer    master_sequencer_D545;
   svt_axi_master_sequencer    master_sequencer_D546;
   svt_axi_master_sequencer    master_sequencer_D547;
   svt_axi_master_sequencer    master_sequencer_D548;
   svt_axi_master_sequencer    master_sequencer_D549;
   svt_axi_master_sequencer    master_sequencer_D550;
   svt_axi_master_sequencer    master_sequencer_D551;
   svt_axi_master_sequencer    master_sequencer_D552;
   svt_axi_master_sequencer    master_sequencer_D553;
   svt_axi_master_sequencer    master_sequencer_D554;
   svt_axi_master_sequencer    master_sequencer_D555;
   svt_axi_master_sequencer    master_sequencer_D556;
   svt_axi_master_sequencer    master_sequencer_D557;
   svt_axi_master_sequencer    master_sequencer_D558;
   svt_axi_master_sequencer    master_sequencer_D559;
   svt_axi_master_sequencer    master_sequencer_D560;
   svt_axi_master_sequencer    master_sequencer_D561;
   svt_axi_master_sequencer    master_sequencer_D562;
   svt_axi_master_sequencer    master_sequencer_D563;
   svt_axi_master_sequencer    master_sequencer_D564;
   svt_axi_master_sequencer    master_sequencer_D565;
   svt_axi_master_sequencer    master_sequencer_D566;
   svt_axi_master_sequencer    master_sequencer_D567;
   svt_axi_master_sequencer    master_sequencer_D568;
   svt_axi_master_sequencer    master_sequencer_D569;
   svt_axi_master_sequencer    master_sequencer_D570;
   svt_axi_master_sequencer    master_sequencer_D571;
   svt_axi_master_sequencer    master_sequencer_D572;
   svt_axi_master_sequencer    master_sequencer_D573;
   svt_axi_master_sequencer    master_sequencer_D574;
   svt_axi_master_sequencer    master_sequencer_D575;
   svt_axi_master_sequencer    master_sequencer_D576;
   svt_axi_master_sequencer    master_sequencer_D577;
   svt_axi_master_sequencer    master_sequencer_D578;
   svt_axi_master_sequencer    master_sequencer_D579;
   svt_axi_master_sequencer    master_sequencer_D580;
   svt_axi_master_sequencer    master_sequencer_D581;
   svt_axi_master_sequencer    master_sequencer_D582;
   svt_axi_master_sequencer    master_sequencer_D583;
   svt_axi_master_sequencer    master_sequencer_D584;
   svt_axi_master_sequencer    master_sequencer_D585;
   svt_axi_master_sequencer    master_sequencer_D586;
   svt_axi_master_sequencer    master_sequencer_D587;
   svt_axi_master_sequencer    master_sequencer_D588;
   svt_axi_master_sequencer    master_sequencer_D589;
   svt_axi_master_sequencer    master_sequencer_D590;
   svt_axi_master_sequencer    master_sequencer_D591;
   svt_axi_master_sequencer    master_sequencer_D592;
   svt_axi_master_sequencer    master_sequencer_D593;
   svt_axi_master_sequencer    master_sequencer_D594;
   svt_axi_master_sequencer    master_sequencer_D595;
   svt_axi_master_sequencer    master_sequencer_D596;
   svt_axi_master_sequencer    master_sequencer_D597;
   svt_axi_master_sequencer    master_sequencer_D598;
   svt_axi_master_sequencer    master_sequencer_D599;
   svt_axi_master_sequencer    master_sequencer_D600;
   svt_axi_master_sequencer    master_sequencer_D601;
   svt_axi_master_sequencer    master_sequencer_D602;
   svt_axi_master_sequencer    master_sequencer_D603;
   svt_axi_master_sequencer    master_sequencer_D604;
   svt_axi_master_sequencer    master_sequencer_D605;
   svt_axi_master_sequencer    master_sequencer_D606;
   svt_axi_master_sequencer    master_sequencer_D607;
   svt_axi_master_sequencer    master_sequencer_D608;
   svt_axi_master_sequencer    master_sequencer_D609;
   svt_axi_master_sequencer    master_sequencer_D610;
   svt_axi_master_sequencer    master_sequencer_D611;
   svt_axi_master_sequencer    master_sequencer_D612;
   svt_axi_master_sequencer    master_sequencer_D613;
   svt_axi_master_sequencer    master_sequencer_D614;
   svt_axi_master_sequencer    master_sequencer_D615;
   svt_axi_master_sequencer    master_sequencer_D616;
   svt_axi_master_sequencer    master_sequencer_D617;
   svt_axi_master_sequencer    master_sequencer_D618;
   svt_axi_master_sequencer    master_sequencer_D619;
   svt_axi_master_sequencer    master_sequencer_D620;
   svt_axi_master_sequencer    master_sequencer_D621;
   svt_axi_master_sequencer    master_sequencer_D622;
   svt_axi_master_sequencer    master_sequencer_D623;
   svt_axi_master_sequencer    master_sequencer_D624;
   svt_axi_master_sequencer    master_sequencer_D625;
   svt_axi_master_sequencer    master_sequencer_D626;
   svt_axi_master_sequencer    master_sequencer_D627;
   svt_axi_master_sequencer    master_sequencer_D628;
   svt_axi_master_sequencer    master_sequencer_D629;
   svt_axi_master_sequencer    master_sequencer_D630;
   svt_axi_master_sequencer    master_sequencer_D631;
   svt_axi_master_sequencer    master_sequencer_D632;
   svt_axi_master_sequencer    master_sequencer_D633;
   svt_axi_master_sequencer    master_sequencer_D634;
   svt_axi_master_sequencer    master_sequencer_D635;
   svt_axi_master_sequencer    master_sequencer_D636;
   svt_axi_master_sequencer    master_sequencer_D637;
   svt_axi_master_sequencer    master_sequencer_D638;
   svt_axi_master_sequencer    master_sequencer_D639;
   svt_axi_master_sequencer    master_sequencer_D640;
   svt_axi_master_sequencer    master_sequencer_D641;
   svt_axi_master_sequencer    master_sequencer_D642;
   svt_axi_master_sequencer    master_sequencer_D643;
   svt_axi_master_sequencer    master_sequencer_D644;
   svt_axi_master_sequencer    master_sequencer_D645;
   svt_axi_master_sequencer    master_sequencer_D646;
   svt_axi_master_sequencer    master_sequencer_D647;
   svt_axi_master_sequencer    master_sequencer_D648;
   svt_axi_master_sequencer    master_sequencer_D649;
   svt_axi_master_sequencer    master_sequencer_D650;
   svt_axi_master_sequencer    master_sequencer_D651;
   svt_axi_master_sequencer    master_sequencer_D652;
   svt_axi_master_sequencer    master_sequencer_D653;
   svt_axi_master_sequencer    master_sequencer_D654;
   svt_axi_master_sequencer    master_sequencer_D655;
   svt_axi_master_sequencer    master_sequencer_D656;
   svt_axi_master_sequencer    master_sequencer_D657;
   svt_axi_master_sequencer    master_sequencer_D658;
   svt_axi_master_sequencer    master_sequencer_D659;
   svt_axi_master_sequencer    master_sequencer_D660;
   svt_axi_master_sequencer    master_sequencer_D661;
   svt_axi_master_sequencer    master_sequencer_D662;
   svt_axi_master_sequencer    master_sequencer_D663;
   svt_axi_master_sequencer    master_sequencer_D664;
   svt_axi_master_sequencer    master_sequencer_D665;
   svt_axi_master_sequencer    master_sequencer_D666;
   svt_axi_master_sequencer    master_sequencer_D667;
   svt_axi_master_sequencer    master_sequencer_D668;
   svt_axi_master_sequencer    master_sequencer_D669;
   svt_axi_master_sequencer    master_sequencer_D670;
   svt_axi_master_sequencer    master_sequencer_D671;
   svt_axi_master_sequencer    master_sequencer_D672;
   svt_axi_master_sequencer    master_sequencer_D673;
   svt_axi_master_sequencer    master_sequencer_D674;
   svt_axi_master_sequencer    master_sequencer_D675;
   svt_axi_master_sequencer    master_sequencer_D676;
   svt_axi_master_sequencer    master_sequencer_D677;
   svt_axi_master_sequencer    master_sequencer_D678;
   svt_axi_master_sequencer    master_sequencer_D679;
   svt_axi_master_sequencer    master_sequencer_D680;
   svt_axi_master_sequencer    master_sequencer_D681;
   svt_axi_master_sequencer    master_sequencer_D682;
   svt_axi_master_sequencer    master_sequencer_D683;
   svt_axi_master_sequencer    master_sequencer_D684;
   svt_axi_master_sequencer    master_sequencer_D685;
   svt_axi_master_sequencer    master_sequencer_D686;
   svt_axi_master_sequencer    master_sequencer_D687;
   svt_axi_master_sequencer    master_sequencer_D688;
   svt_axi_master_sequencer    master_sequencer_D689;
   svt_axi_master_sequencer    master_sequencer_D690;
   svt_axi_master_sequencer    master_sequencer_D691;
   svt_axi_master_sequencer    master_sequencer_D692;
   svt_axi_master_sequencer    master_sequencer_D693;
   svt_axi_master_sequencer    master_sequencer_D694;
   svt_axi_master_sequencer    master_sequencer_D695;
   svt_axi_master_sequencer    master_sequencer_D696;
   svt_axi_master_sequencer    master_sequencer_D697;
   svt_axi_master_sequencer    master_sequencer_D698;
   svt_axi_master_sequencer    master_sequencer_D699;
   svt_axi_master_sequencer    master_sequencer_D700;
   svt_axi_master_sequencer    master_sequencer_D701;
   svt_axi_master_sequencer    master_sequencer_D702;
   svt_axi_master_sequencer    master_sequencer_D703;
   svt_axi_master_sequencer    master_sequencer_D704;
   svt_axi_master_sequencer    master_sequencer_D705;
   svt_axi_master_sequencer    master_sequencer_D706;
   svt_axi_master_sequencer    master_sequencer_D707;
   svt_axi_master_sequencer    master_sequencer_D708;
   svt_axi_master_sequencer    master_sequencer_D709;
   svt_axi_master_sequencer    master_sequencer_D710;
   svt_axi_master_sequencer    master_sequencer_D711;
   svt_axi_master_sequencer    master_sequencer_D712;
   svt_axi_master_sequencer    master_sequencer_D713;
   svt_axi_master_sequencer    master_sequencer_D714;
   svt_axi_master_sequencer    master_sequencer_D715;
   svt_axi_master_sequencer    master_sequencer_D716;
   svt_axi_master_sequencer    master_sequencer_D717;
   svt_axi_master_sequencer    master_sequencer_D718;
   svt_axi_master_sequencer    master_sequencer_D719;
   svt_axi_master_sequencer    master_sequencer_D720;
   svt_axi_master_sequencer    master_sequencer_D721;
   svt_axi_master_sequencer    master_sequencer_D722;
   svt_axi_master_sequencer    master_sequencer_D723;
   svt_axi_master_sequencer    master_sequencer_D724;
   svt_axi_master_sequencer    master_sequencer_D725;
   svt_axi_master_sequencer    master_sequencer_D726;
   svt_axi_master_sequencer    master_sequencer_D727;
   svt_axi_master_sequencer    master_sequencer_D728;
   svt_axi_master_sequencer    master_sequencer_D729;
   svt_axi_master_sequencer    master_sequencer_D730;
   svt_axi_master_sequencer    master_sequencer_D731;
   svt_axi_master_sequencer    master_sequencer_D732;
   svt_axi_master_sequencer    master_sequencer_D733;
   svt_axi_master_sequencer    master_sequencer_D734;
   svt_axi_master_sequencer    master_sequencer_D735;
   svt_axi_master_sequencer    master_sequencer_D736;
   svt_axi_master_sequencer    master_sequencer_D737;
   svt_axi_master_sequencer    master_sequencer_D738;
   svt_axi_master_sequencer    master_sequencer_D739;
   svt_axi_master_sequencer    master_sequencer_D740;
   svt_axi_master_sequencer    master_sequencer_D741;
   svt_axi_master_sequencer    master_sequencer_D742;
   svt_axi_master_sequencer    master_sequencer_D743;
   svt_axi_master_sequencer    master_sequencer_D744;
   svt_axi_master_sequencer    master_sequencer_D745;
   svt_axi_master_sequencer    master_sequencer_D746;
   svt_axi_master_sequencer    master_sequencer_D747;
   svt_axi_master_sequencer    master_sequencer_D748;
   svt_axi_master_sequencer    master_sequencer_D749;
   svt_axi_master_sequencer    master_sequencer_D750;
   svt_axi_master_sequencer    master_sequencer_D751;
   svt_axi_master_sequencer    master_sequencer_D752;
   svt_axi_master_sequencer    master_sequencer_D753;
   svt_axi_master_sequencer    master_sequencer_D754;
   svt_axi_master_sequencer    master_sequencer_D755;
   svt_axi_master_sequencer    master_sequencer_D756;
   svt_axi_master_sequencer    master_sequencer_D757;
   svt_axi_master_sequencer    master_sequencer_D758;
   svt_axi_master_sequencer    master_sequencer_D759;
   svt_axi_master_sequencer    master_sequencer_D760;
   svt_axi_master_sequencer    master_sequencer_D761;
   svt_axi_master_sequencer    master_sequencer_D762;
   svt_axi_master_sequencer    master_sequencer_D763;
   svt_axi_master_sequencer    master_sequencer_D764;
   svt_axi_master_sequencer    master_sequencer_D765;
   svt_axi_master_sequencer    master_sequencer_D766;
   svt_axi_master_sequencer    master_sequencer_D767;
   svt_axi_master_sequencer    master_sequencer_D768;
   svt_axi_master_sequencer    master_sequencer_D769;
   svt_axi_master_sequencer    master_sequencer_D770;
   svt_axi_master_sequencer    master_sequencer_D771;
   svt_axi_master_sequencer    master_sequencer_D772;
   svt_axi_master_sequencer    master_sequencer_D773;
   svt_axi_master_sequencer    master_sequencer_D774;
   svt_axi_master_sequencer    master_sequencer_D775;
   svt_axi_master_sequencer    master_sequencer_D776;
   svt_axi_master_sequencer    master_sequencer_D777;
   svt_axi_master_sequencer    master_sequencer_D778;
   svt_axi_master_sequencer    master_sequencer_D779;
   svt_axi_master_sequencer    master_sequencer_D780;
   svt_axi_master_sequencer    master_sequencer_D781;
   svt_axi_master_sequencer    master_sequencer_D782;
   svt_axi_master_sequencer    master_sequencer_D783;
   svt_axi_master_sequencer    master_sequencer_D784;
   svt_axi_master_sequencer    master_sequencer_D785;
   svt_axi_master_sequencer    master_sequencer_D786;
   svt_axi_master_sequencer    master_sequencer_D787;
   svt_axi_master_sequencer    master_sequencer_D788;
   svt_axi_master_sequencer    master_sequencer_D789;
   svt_axi_master_sequencer    master_sequencer_D790;
   svt_axi_master_sequencer    master_sequencer_D791;
   svt_axi_master_sequencer    master_sequencer_D792;
   svt_axi_master_sequencer    master_sequencer_D793;
   svt_axi_master_sequencer    master_sequencer_D794;
   svt_axi_master_sequencer    master_sequencer_D795;
   svt_axi_master_sequencer    master_sequencer_D796;
   svt_axi_master_sequencer    master_sequencer_D797;
   svt_axi_master_sequencer    master_sequencer_D798;
   svt_axi_master_sequencer    master_sequencer_D799;
   svt_axi_master_sequencer    master_sequencer_D800;
   svt_axi_master_sequencer    master_sequencer_D801;
   svt_axi_master_sequencer    master_sequencer_D802;
   svt_axi_master_sequencer    master_sequencer_D803;
   svt_axi_master_sequencer    master_sequencer_D804;
   svt_axi_master_sequencer    master_sequencer_D805;
   svt_axi_master_sequencer    master_sequencer_D806;
   svt_axi_master_sequencer    master_sequencer_D807;
   svt_axi_master_sequencer    master_sequencer_D808;
   svt_axi_master_sequencer    master_sequencer_D809;
   svt_axi_master_sequencer    master_sequencer_D810;
   svt_axi_master_sequencer    master_sequencer_D811;
   svt_axi_master_sequencer    master_sequencer_D812;
   svt_axi_master_sequencer    master_sequencer_D813;
   svt_axi_master_sequencer    master_sequencer_D814;
   svt_axi_master_sequencer    master_sequencer_D815;
   svt_axi_master_sequencer    master_sequencer_D816;
   svt_axi_master_sequencer    master_sequencer_D817;
   svt_axi_master_sequencer    master_sequencer_D818;
   svt_axi_master_sequencer    master_sequencer_D819;
   svt_axi_master_sequencer    master_sequencer_D820;
   svt_axi_master_sequencer    master_sequencer_D821;
   svt_axi_master_sequencer    master_sequencer_D822;
   svt_axi_master_sequencer    master_sequencer_D823;
   svt_axi_master_sequencer    master_sequencer_D824;
   svt_axi_master_sequencer    master_sequencer_D825;
   svt_axi_master_sequencer    master_sequencer_D826;
   svt_axi_master_sequencer    master_sequencer_D827;
   svt_axi_master_sequencer    master_sequencer_D828;
   svt_axi_master_sequencer    master_sequencer_D829;
   svt_axi_master_sequencer    master_sequencer_D830;
   svt_axi_master_sequencer    master_sequencer_D831;
   svt_axi_master_sequencer    master_sequencer_D832;
   svt_axi_master_sequencer    master_sequencer_D833;
   svt_axi_master_sequencer    master_sequencer_D834;
   svt_axi_master_sequencer    master_sequencer_D835;
   svt_axi_master_sequencer    master_sequencer_D836;
   svt_axi_master_sequencer    master_sequencer_D837;
   svt_axi_master_sequencer    master_sequencer_D838;
   svt_axi_master_sequencer    master_sequencer_D839;
   svt_axi_master_sequencer    master_sequencer_D840;
   svt_axi_master_sequencer    master_sequencer_D841;
   svt_axi_master_sequencer    master_sequencer_D842;
   svt_axi_master_sequencer    master_sequencer_D843;
   svt_axi_master_sequencer    master_sequencer_D844;
   svt_axi_master_sequencer    master_sequencer_D845;
   svt_axi_master_sequencer    master_sequencer_D846;
   svt_axi_master_sequencer    master_sequencer_D847;
   svt_axi_master_sequencer    master_sequencer_D848;
   svt_axi_master_sequencer    master_sequencer_D849;
   svt_axi_master_sequencer    master_sequencer_D850;
   svt_axi_master_sequencer    master_sequencer_D851;
   svt_axi_master_sequencer    master_sequencer_D852;
   svt_axi_master_sequencer    master_sequencer_D853;
   svt_axi_master_sequencer    master_sequencer_D854;
   svt_axi_master_sequencer    master_sequencer_D855;
   svt_axi_master_sequencer    master_sequencer_D856;
   svt_axi_master_sequencer    master_sequencer_D857;
   svt_axi_master_sequencer    master_sequencer_D858;
   svt_axi_master_sequencer    master_sequencer_D859;
   svt_axi_master_sequencer    master_sequencer_D860;
   svt_axi_master_sequencer    master_sequencer_D861;
   svt_axi_master_sequencer    master_sequencer_D862;
   svt_axi_master_sequencer    master_sequencer_D863;
   svt_axi_master_sequencer    master_sequencer_D864;
   svt_axi_master_sequencer    master_sequencer_D865;
   svt_axi_master_sequencer    master_sequencer_D866;
   svt_axi_master_sequencer    master_sequencer_D867;
   svt_axi_master_sequencer    master_sequencer_D868;
   svt_axi_master_sequencer    master_sequencer_D869;
   svt_axi_master_sequencer    master_sequencer_D870;
   svt_axi_master_sequencer    master_sequencer_D871;
   svt_axi_master_sequencer    master_sequencer_D872;
   svt_axi_master_sequencer    master_sequencer_D873;
   svt_axi_master_sequencer    master_sequencer_D874;
   svt_axi_master_sequencer    master_sequencer_D875;
   svt_axi_master_sequencer    master_sequencer_D876;
   svt_axi_master_sequencer    master_sequencer_D877;
   svt_axi_master_sequencer    master_sequencer_D878;
   svt_axi_master_sequencer    master_sequencer_D879;
   svt_axi_master_sequencer    master_sequencer_D880;
   svt_axi_master_sequencer    master_sequencer_D881;
   svt_axi_master_sequencer    master_sequencer_D882;
   svt_axi_master_sequencer    master_sequencer_D883;
   svt_axi_master_sequencer    master_sequencer_D884;
   svt_axi_master_sequencer    master_sequencer_D885;
   svt_axi_master_sequencer    master_sequencer_D886;
   svt_axi_master_sequencer    master_sequencer_D887;
   svt_axi_master_sequencer    master_sequencer_D888;
   svt_axi_master_sequencer    master_sequencer_D889;
   svt_axi_master_sequencer    master_sequencer_D890;
   svt_axi_master_sequencer    master_sequencer_D891;
   svt_axi_master_sequencer    master_sequencer_D892;
   svt_axi_master_sequencer    master_sequencer_D893;
   svt_axi_master_sequencer    master_sequencer_D894;
   svt_axi_master_sequencer    master_sequencer_D895;
   svt_axi_master_sequencer    master_sequencer_D896;
   svt_axi_master_sequencer    master_sequencer_D897;
   svt_axi_master_sequencer    master_sequencer_D898;
   svt_axi_master_sequencer    master_sequencer_D899;
   svt_axi_master_sequencer    master_sequencer_D900;
   svt_axi_master_sequencer    master_sequencer_D901;
   svt_axi_master_sequencer    master_sequencer_D902;
   svt_axi_master_sequencer    master_sequencer_D903;
   svt_axi_master_sequencer    master_sequencer_D904;
   svt_axi_master_sequencer    master_sequencer_D905;
   svt_axi_master_sequencer    master_sequencer_D906;
   svt_axi_master_sequencer    master_sequencer_D907;
   svt_axi_master_sequencer    master_sequencer_D908;
   svt_axi_master_sequencer    master_sequencer_D909;
   svt_axi_master_sequencer    master_sequencer_D910;
   svt_axi_master_sequencer    master_sequencer_D911;
   svt_axi_master_sequencer    master_sequencer_D912;
   svt_axi_master_sequencer    master_sequencer_D913;
   svt_axi_master_sequencer    master_sequencer_D914;
   svt_axi_master_sequencer    master_sequencer_D915;
   svt_axi_master_sequencer    master_sequencer_D916;
   svt_axi_master_sequencer    master_sequencer_D917;
   svt_axi_master_sequencer    master_sequencer_D918;
   svt_axi_master_sequencer    master_sequencer_D919;
   svt_axi_master_sequencer    master_sequencer_D920;
   svt_axi_master_sequencer    master_sequencer_D921;
   svt_axi_master_sequencer    master_sequencer_D922;
   svt_axi_master_sequencer    master_sequencer_D923;
   svt_axi_master_sequencer    master_sequencer_D924;
   svt_axi_master_sequencer    master_sequencer_D925;
   svt_axi_master_sequencer    master_sequencer_D926;
   svt_axi_master_sequencer    master_sequencer_D927;
   svt_axi_master_sequencer    master_sequencer_D928;
   svt_axi_master_sequencer    master_sequencer_D929;
   svt_axi_master_sequencer    master_sequencer_D930;
   svt_axi_master_sequencer    master_sequencer_D931;
   svt_axi_master_sequencer    master_sequencer_D932;
   svt_axi_master_sequencer    master_sequencer_D933;
   svt_axi_master_sequencer    master_sequencer_D934;
   svt_axi_master_sequencer    master_sequencer_D935;
   svt_axi_master_sequencer    master_sequencer_D936;
   svt_axi_master_sequencer    master_sequencer_D937;
   svt_axi_master_sequencer    master_sequencer_D938;
   svt_axi_master_sequencer    master_sequencer_D939;
   svt_axi_master_sequencer    master_sequencer_D940;
   svt_axi_master_sequencer    master_sequencer_D941;
   svt_axi_master_sequencer    master_sequencer_D942;
   svt_axi_master_sequencer    master_sequencer_D943;
   svt_axi_master_sequencer    master_sequencer_D944;
   svt_axi_master_sequencer    master_sequencer_D945;
   svt_axi_master_sequencer    master_sequencer_D946;
   svt_axi_master_sequencer    master_sequencer_D947;
   svt_axi_master_sequencer    master_sequencer_D948;
   svt_axi_master_sequencer    master_sequencer_D949;
   svt_axi_master_sequencer    master_sequencer_D950;
   svt_axi_master_sequencer    master_sequencer_D951;
   svt_axi_master_sequencer    master_sequencer_D952;
   svt_axi_master_sequencer    master_sequencer_D953;
   svt_axi_master_sequencer    master_sequencer_D954;
   svt_axi_master_sequencer    master_sequencer_D955;
   svt_axi_master_sequencer    master_sequencer_D956;
   svt_axi_master_sequencer    master_sequencer_D957;
   svt_axi_master_sequencer    master_sequencer_D958;
   svt_axi_master_sequencer    master_sequencer_D959;
   svt_axi_master_sequencer    master_sequencer_D960;
   svt_axi_master_sequencer    master_sequencer_D961;
   svt_axi_master_sequencer    master_sequencer_D962;
   svt_axi_master_sequencer    master_sequencer_D963;
   svt_axi_master_sequencer    master_sequencer_D964;
   svt_axi_master_sequencer    master_sequencer_D965;
   svt_axi_master_sequencer    master_sequencer_D966;
   svt_axi_master_sequencer    master_sequencer_D967;
   svt_axi_master_sequencer    master_sequencer_D968;
   svt_axi_master_sequencer    master_sequencer_D969;
   svt_axi_master_sequencer    master_sequencer_D970;
   svt_axi_master_sequencer    master_sequencer_D971;
   svt_axi_master_sequencer    master_sequencer_D972;
   svt_axi_master_sequencer    master_sequencer_D973;
   svt_axi_master_sequencer    master_sequencer_D974;
   svt_axi_master_sequencer    master_sequencer_D975;
   svt_axi_master_sequencer    master_sequencer_D976;
   svt_axi_master_sequencer    master_sequencer_D977;
   svt_axi_master_sequencer    master_sequencer_D978;
   svt_axi_master_sequencer    master_sequencer_D979;
   svt_axi_master_sequencer    master_sequencer_D980;
   svt_axi_master_sequencer    master_sequencer_D981;
   svt_axi_master_sequencer    master_sequencer_D982;
   svt_axi_master_sequencer    master_sequencer_D983;
   svt_axi_master_sequencer    master_sequencer_D984;
   svt_axi_master_sequencer    master_sequencer_D985;
   svt_axi_master_sequencer    master_sequencer_D986;
   svt_axi_master_sequencer    master_sequencer_D987;
   svt_axi_master_sequencer    master_sequencer_D988;
   svt_axi_master_sequencer    master_sequencer_D989;
   svt_axi_master_sequencer    master_sequencer_D990;
   svt_axi_master_sequencer    master_sequencer_D991;
   svt_axi_master_sequencer    master_sequencer_D992;
   svt_axi_master_sequencer    master_sequencer_D993;
   svt_axi_master_sequencer    master_sequencer_D994;
   svt_axi_master_sequencer    master_sequencer_D995;
   svt_axi_master_sequencer    master_sequencer_D996;
   svt_axi_master_sequencer    master_sequencer_D997;
   svt_axi_master_sequencer    master_sequencer_D998;
   svt_axi_master_sequencer    master_sequencer_D999;
   svt_axi_master_sequencer    master_sequencer_D1000;
   svt_axi_master_sequencer    master_sequencer_D1001;
   svt_axi_master_sequencer    master_sequencer_D1002;
   svt_axi_master_sequencer    master_sequencer_D1003;
   svt_axi_master_sequencer    master_sequencer_D1004;
   svt_axi_master_sequencer    master_sequencer_D1005;
   svt_axi_master_sequencer    master_sequencer_D1006;
   svt_axi_master_sequencer    master_sequencer_D1007;
   svt_axi_master_sequencer    master_sequencer_D1008;
   svt_axi_master_sequencer    master_sequencer_D1009;
   svt_axi_master_sequencer    master_sequencer_D1010;
   svt_axi_master_sequencer    master_sequencer_D1011;
   svt_axi_master_sequencer    master_sequencer_D1012;
   svt_axi_master_sequencer    master_sequencer_D1013;
   svt_axi_master_sequencer    master_sequencer_D1014;
   svt_axi_master_sequencer    master_sequencer_D1015;
   svt_axi_master_sequencer    master_sequencer_D1016;
   svt_axi_master_sequencer    master_sequencer_D1017;
   svt_axi_master_sequencer    master_sequencer_D1018;
   svt_axi_master_sequencer    master_sequencer_D1019;
   svt_axi_master_sequencer    master_sequencer_D1020;
   svt_axi_master_sequencer    master_sequencer_D1021;
   svt_axi_master_sequencer    master_sequencer_D1022;
   svt_axi_master_sequencer    master_sequencer_D1023;
   svt_axi_master_sequencer    master_sequencer_D1024;
   svt_axi_master_sequencer    master_sequencer_D1025;
   svt_axi_master_sequencer    master_sequencer_D1026;
   svt_axi_master_sequencer    master_sequencer_D1027;
   svt_axi_master_sequencer    master_sequencer_D1028;
   svt_axi_master_sequencer    master_sequencer_D1029;
   svt_axi_master_sequencer    master_sequencer_D1030;
   svt_axi_master_sequencer    master_sequencer_D1031;
   svt_axi_master_sequencer    master_sequencer_D1032;
   svt_axi_master_sequencer    master_sequencer_D1033;
   svt_axi_master_sequencer    master_sequencer_D1034;
   svt_axi_master_sequencer    master_sequencer_D1035;
   svt_axi_master_sequencer    master_sequencer_D1036;
   svt_axi_master_sequencer    master_sequencer_D1037;
   svt_axi_master_sequencer    master_sequencer_D1038;
   svt_axi_master_sequencer    master_sequencer_D1039;
   svt_axi_master_sequencer    master_sequencer_D1040;
   svt_axi_master_sequencer    master_sequencer_D1041;
   svt_axi_master_sequencer    master_sequencer_D1042;
   svt_axi_master_sequencer    master_sequencer_D1043;
   svt_axi_master_sequencer    master_sequencer_D1044;
   svt_axi_master_sequencer    master_sequencer_D1045;
   svt_axi_master_sequencer    master_sequencer_D1046;
   svt_axi_master_sequencer    master_sequencer_D1047;
   svt_axi_master_sequencer    master_sequencer_D1048;
   svt_axi_master_sequencer    master_sequencer_D1049;
   svt_axi_master_sequencer    master_sequencer_D1050;
   svt_axi_master_sequencer    master_sequencer_D1051;
   svt_axi_master_sequencer    master_sequencer_D1052;
   svt_axi_master_sequencer    master_sequencer_D1053;
   svt_axi_master_sequencer    master_sequencer_D1054;
   svt_axi_master_sequencer    master_sequencer_D1055;
   svt_axi_master_sequencer    master_sequencer_D1056;
   svt_axi_master_sequencer    master_sequencer_D1057;
   svt_axi_master_sequencer    master_sequencer_D1058;
   svt_axi_master_sequencer    master_sequencer_D1059;
   svt_axi_master_sequencer    master_sequencer_D1060;
   svt_axi_master_sequencer    master_sequencer_D1061;
   svt_axi_master_sequencer    master_sequencer_D1062;
   svt_axi_master_sequencer    master_sequencer_D1063;
   svt_axi_master_sequencer    master_sequencer_D1064;
   svt_axi_master_sequencer    master_sequencer_D1065;
   svt_axi_master_sequencer    master_sequencer_D1066;
   svt_axi_master_sequencer    master_sequencer_D1067;
   svt_axi_master_sequencer    master_sequencer_D1068;
   svt_axi_master_sequencer    master_sequencer_D1069;
   svt_axi_master_sequencer    master_sequencer_D1070;
   svt_axi_master_sequencer    master_sequencer_D1071;
   svt_axi_master_sequencer    master_sequencer_D1072;
   svt_axi_master_sequencer    master_sequencer_D1073;
   svt_axi_master_sequencer    master_sequencer_D1074;
   svt_axi_master_sequencer    master_sequencer_D1075;
   svt_axi_master_sequencer    master_sequencer_D1076;
   svt_axi_master_sequencer    master_sequencer_D1077;
   svt_axi_master_sequencer    master_sequencer_D1078;
   svt_axi_master_sequencer    master_sequencer_D1079;
   svt_axi_master_sequencer    master_sequencer_D1080;
   svt_axi_master_sequencer    master_sequencer_D1081;
   svt_axi_master_sequencer    master_sequencer_D1082;
   svt_axi_master_sequencer    master_sequencer_D1083;
   svt_axi_master_sequencer    master_sequencer_D1084;
   svt_axi_master_sequencer    master_sequencer_D1085;
   svt_axi_master_sequencer    master_sequencer_D1086;
   svt_axi_master_sequencer    master_sequencer_D1087;
   svt_axi_master_sequencer    master_sequencer_D1088;
   svt_axi_master_sequencer    master_sequencer_D1089;
   svt_axi_master_sequencer    master_sequencer_D1090;
   svt_axi_master_sequencer    master_sequencer_D1091;
   svt_axi_master_sequencer    master_sequencer_D1092;
   svt_axi_master_sequencer    master_sequencer_D1093;
   svt_axi_master_sequencer    master_sequencer_D1094;
   svt_axi_master_sequencer    master_sequencer_D1095;
   svt_axi_master_sequencer    master_sequencer_D1096;
   svt_axi_master_sequencer    master_sequencer_D1097;
   svt_axi_master_sequencer    master_sequencer_D1098;
   svt_axi_master_sequencer    master_sequencer_D1099;
   svt_axi_master_sequencer    master_sequencer_D1100;
   svt_axi_master_sequencer    master_sequencer_D1101;
   svt_axi_master_sequencer    master_sequencer_D1102;
   svt_axi_master_sequencer    master_sequencer_D1103;
   svt_axi_master_sequencer    master_sequencer_D1104;
   svt_axi_master_sequencer    master_sequencer_D1105;
   svt_axi_master_sequencer    master_sequencer_D1106;
   svt_axi_master_sequencer    master_sequencer_D1107;
   svt_axi_master_sequencer    master_sequencer_D1108;
   svt_axi_master_sequencer    master_sequencer_D1109;
   svt_axi_master_sequencer    master_sequencer_D1110;
   svt_axi_master_sequencer    master_sequencer_D1111;
   svt_axi_master_sequencer    master_sequencer_D1112;
   svt_axi_master_sequencer    master_sequencer_D1113;
   svt_axi_master_sequencer    master_sequencer_D1114;
   svt_axi_master_sequencer    master_sequencer_D1115;
   svt_axi_master_sequencer    master_sequencer_D1116;
   svt_axi_master_sequencer    master_sequencer_D1117;
   svt_axi_master_sequencer    master_sequencer_D1118;
   svt_axi_master_sequencer    master_sequencer_D1119;
   svt_axi_master_sequencer    master_sequencer_D1120;
   svt_axi_master_sequencer    master_sequencer_D1121;
   svt_axi_master_sequencer    master_sequencer_D1122;
   svt_axi_master_sequencer    master_sequencer_D1123;
   svt_axi_master_sequencer    master_sequencer_D1124;
   svt_axi_master_sequencer    master_sequencer_D1125;
   svt_axi_master_sequencer    master_sequencer_D1126;
   svt_axi_master_sequencer    master_sequencer_D1127;
   svt_axi_master_sequencer    master_sequencer_D1128;
   svt_axi_master_sequencer    master_sequencer_D1129;
   svt_axi_master_sequencer    master_sequencer_D1130;
   svt_axi_master_sequencer    master_sequencer_D1131;
   svt_axi_master_sequencer    master_sequencer_D1132;
   svt_axi_master_sequencer    master_sequencer_D1133;
   svt_axi_master_sequencer    master_sequencer_D1134;
   svt_axi_master_sequencer    master_sequencer_D1135;
   svt_axi_master_sequencer    master_sequencer_D1136;
   svt_axi_master_sequencer    master_sequencer_D1137;
   svt_axi_master_sequencer    master_sequencer_D1138;
   svt_axi_master_sequencer    master_sequencer_D1139;
   svt_axi_master_sequencer    master_sequencer_D1140;
   svt_axi_master_sequencer    master_sequencer_D1141;
   svt_axi_master_sequencer    master_sequencer_D1142;
   svt_axi_master_sequencer    master_sequencer_D1143;
   svt_axi_master_sequencer    master_sequencer_D1144;
   svt_axi_master_sequencer    master_sequencer_D1145;
   svt_axi_master_sequencer    master_sequencer_D1146;
   svt_axi_master_sequencer    master_sequencer_D1147;
   svt_axi_master_sequencer    master_sequencer_D1148;
   svt_axi_master_sequencer    master_sequencer_D1149;
   svt_axi_master_sequencer    master_sequencer_D1150;
   svt_axi_master_sequencer    master_sequencer_D1151;
   svt_axi_master_sequencer    master_sequencer_D1152;
   svt_axi_master_sequencer    master_sequencer_D1153;
   svt_axi_master_sequencer    master_sequencer_D1154;
   svt_axi_master_sequencer    master_sequencer_D1155;
   svt_axi_master_sequencer    master_sequencer_D1156;
   svt_axi_master_sequencer    master_sequencer_D1157;
   svt_axi_master_sequencer    master_sequencer_D1158;
   svt_axi_master_sequencer    master_sequencer_D1159;
   svt_axi_master_sequencer    master_sequencer_D1160;
   svt_axi_master_sequencer    master_sequencer_D1161;
   svt_axi_master_sequencer    master_sequencer_D1162;
   svt_axi_master_sequencer    master_sequencer_D1163;
   svt_axi_master_sequencer    master_sequencer_D1164;
   svt_axi_master_sequencer    master_sequencer_D1165;
   svt_axi_master_sequencer    master_sequencer_D1166;
   svt_axi_master_sequencer    master_sequencer_D1167;
   svt_axi_master_sequencer    master_sequencer_D1168;
   svt_axi_master_sequencer    master_sequencer_D1169;
   svt_axi_master_sequencer    master_sequencer_D1170;
   svt_axi_master_sequencer    master_sequencer_D1171;
   svt_axi_master_sequencer    master_sequencer_D1172;
   svt_axi_master_sequencer    master_sequencer_D1173;
   svt_axi_master_sequencer    master_sequencer_D1174;
   svt_axi_master_sequencer    master_sequencer_D1175;
   svt_axi_master_sequencer    master_sequencer_D1176;
   svt_axi_master_sequencer    master_sequencer_D1177;
   svt_axi_master_sequencer    master_sequencer_D1178;
   svt_axi_master_sequencer    master_sequencer_D1179;
   svt_axi_master_sequencer    master_sequencer_D1180;
   svt_axi_master_sequencer    master_sequencer_D1181;
   svt_axi_master_sequencer    master_sequencer_D1182;
   svt_axi_master_sequencer    master_sequencer_D1183;
   svt_axi_master_sequencer    master_sequencer_D1184;
   svt_axi_master_sequencer    master_sequencer_D1185;
   svt_axi_master_sequencer    master_sequencer_D1186;
   svt_axi_master_sequencer    master_sequencer_D1187;
   svt_axi_master_sequencer    master_sequencer_D1188;
   svt_axi_master_sequencer    master_sequencer_D1189;
   svt_axi_master_sequencer    master_sequencer_D1190;
   svt_axi_master_sequencer    master_sequencer_D1191;
   svt_axi_master_sequencer    master_sequencer_D1192;
   svt_axi_master_sequencer    master_sequencer_D1193;
   svt_axi_master_sequencer    master_sequencer_D1194;
   svt_axi_master_sequencer    master_sequencer_D1195;
   svt_axi_master_sequencer    master_sequencer_D1196;
   svt_axi_master_sequencer    master_sequencer_D1197;
   svt_axi_master_sequencer    master_sequencer_D1198;
   svt_axi_master_sequencer    master_sequencer_D1199;
   svt_axi_master_sequencer    master_sequencer_D1200;
   svt_axi_master_sequencer    master_sequencer_D1201;
   svt_axi_master_sequencer    master_sequencer_D1202;
   svt_axi_master_sequencer    master_sequencer_D1203;
   svt_axi_master_sequencer    master_sequencer_D1204;
   svt_axi_master_sequencer    master_sequencer_D1205;
   svt_axi_master_sequencer    master_sequencer_D1206;
   svt_axi_master_sequencer    master_sequencer_D1207;
   svt_axi_master_sequencer    master_sequencer_D1208;
   svt_axi_master_sequencer    master_sequencer_D1209;
   svt_axi_master_sequencer    master_sequencer_D1210;
   svt_axi_master_sequencer    master_sequencer_D1211;
   svt_axi_master_sequencer    master_sequencer_D1212;
   svt_axi_master_sequencer    master_sequencer_D1213;
   svt_axi_master_sequencer    master_sequencer_D1214;
   svt_axi_master_sequencer    master_sequencer_D1215;
   svt_axi_master_sequencer    master_sequencer_D1216;
   svt_axi_master_sequencer    master_sequencer_D1217;
   svt_axi_master_sequencer    master_sequencer_D1218;
   svt_axi_master_sequencer    master_sequencer_D1219;
   svt_axi_master_sequencer    master_sequencer_D1220;
   svt_axi_master_sequencer    master_sequencer_D1221;
   svt_axi_master_sequencer    master_sequencer_D1222;
   svt_axi_master_sequencer    master_sequencer_D1223;
   svt_axi_master_sequencer    master_sequencer_D1224;
   svt_axi_master_sequencer    master_sequencer_D1225;
   svt_axi_master_sequencer    master_sequencer_D1226;
   svt_axi_master_sequencer    master_sequencer_D1227;
   svt_axi_master_sequencer    master_sequencer_D1228;
   svt_axi_master_sequencer    master_sequencer_D1229;
   svt_axi_master_sequencer    master_sequencer_D1230;
   svt_axi_master_sequencer    master_sequencer_D1231;
   svt_axi_master_sequencer    master_sequencer_D1232;
   svt_axi_master_sequencer    master_sequencer_D1233;
   svt_axi_master_sequencer    master_sequencer_D1234;
   svt_axi_master_sequencer    master_sequencer_D1235;
   svt_axi_master_sequencer    master_sequencer_D1236;
   svt_axi_master_sequencer    master_sequencer_D1237;
   svt_axi_master_sequencer    master_sequencer_D1238;
   svt_axi_master_sequencer    master_sequencer_D1239;
   svt_axi_master_sequencer    master_sequencer_D1240;
   svt_axi_master_sequencer    master_sequencer_D1241;
   svt_axi_master_sequencer    master_sequencer_D1242;
   svt_axi_master_sequencer    master_sequencer_D1243;
   svt_axi_master_sequencer    master_sequencer_D1244;
   svt_axi_master_sequencer    master_sequencer_D1245;
   svt_axi_master_sequencer    master_sequencer_D1246;
   svt_axi_master_sequencer    master_sequencer_D1247;
   svt_axi_master_sequencer    master_sequencer_D1248;
   svt_axi_master_sequencer    master_sequencer_D1249;
   svt_axi_master_sequencer    master_sequencer_D1250;
   svt_axi_master_sequencer    master_sequencer_D1251;
   svt_axi_master_sequencer    master_sequencer_D1252;
   svt_axi_master_sequencer    master_sequencer_D1253;
   svt_axi_master_sequencer    master_sequencer_D1254;
   svt_axi_master_sequencer    master_sequencer_D1255;
   svt_axi_master_sequencer    master_sequencer_D1256;
   svt_axi_master_sequencer    master_sequencer_D1257;
   svt_axi_master_sequencer    master_sequencer_D1258;
   svt_axi_master_sequencer    master_sequencer_D1259;
   svt_axi_master_sequencer    master_sequencer_D1260;
   svt_axi_master_sequencer    master_sequencer_D1261;
   svt_axi_master_sequencer    master_sequencer_D1262;
   svt_axi_master_sequencer    master_sequencer_D1263;
   svt_axi_master_sequencer    master_sequencer_D1264;
   svt_axi_master_sequencer    master_sequencer_D1265;
   svt_axi_master_sequencer    master_sequencer_D1266;
   svt_axi_master_sequencer    master_sequencer_D1267;
   svt_axi_master_sequencer    master_sequencer_D1268;
   svt_axi_master_sequencer    master_sequencer_D1269;
   svt_axi_master_sequencer    master_sequencer_D1270;
   svt_axi_master_sequencer    master_sequencer_D1271;
   svt_axi_master_sequencer    master_sequencer_D1272;
   svt_axi_master_sequencer    master_sequencer_D1273;
   svt_axi_master_sequencer    master_sequencer_D1274;
   svt_axi_master_sequencer    master_sequencer_D1275;
   svt_axi_master_sequencer    master_sequencer_D1276;
   svt_axi_master_sequencer    master_sequencer_D1277;
   svt_axi_master_sequencer    master_sequencer_D1278;
   svt_axi_master_sequencer    master_sequencer_D1279;
   svt_axi_master_sequencer    master_sequencer_D1280;
   svt_axi_master_sequencer    master_sequencer_D1281;
   svt_axi_master_sequencer    master_sequencer_D1282;
   svt_axi_master_sequencer    master_sequencer_D1283;
   svt_axi_master_sequencer    master_sequencer_D1284;
   svt_axi_master_sequencer    master_sequencer_D1285;
   svt_axi_master_sequencer    master_sequencer_D1286;
   svt_axi_master_sequencer    master_sequencer_D1287;
   svt_axi_master_sequencer    master_sequencer_D1288;
   svt_axi_master_sequencer    master_sequencer_D1289;
   svt_axi_master_sequencer    master_sequencer_D1290;
   svt_axi_master_sequencer    master_sequencer_D1291;
   svt_axi_master_sequencer    master_sequencer_D1292;
   svt_axi_master_sequencer    master_sequencer_D1293;
   svt_axi_master_sequencer    master_sequencer_D1294;
   svt_axi_master_sequencer    master_sequencer_D1295;
   svt_axi_master_sequencer    master_sequencer_D1296;
   svt_axi_master_sequencer    master_sequencer_D1297;
   svt_axi_master_sequencer    master_sequencer_D1298;
   svt_axi_master_sequencer    master_sequencer_D1299;
   svt_axi_master_sequencer    master_sequencer_D1300;
   svt_axi_master_sequencer    master_sequencer_D1301;
   svt_axi_master_sequencer    master_sequencer_D1302;
   svt_axi_master_sequencer    master_sequencer_D1303;
   svt_axi_master_sequencer    master_sequencer_D1304;
   svt_axi_master_sequencer    master_sequencer_D1305;
   svt_axi_master_sequencer    master_sequencer_D1306;
   svt_axi_master_sequencer    master_sequencer_D1307;
   svt_axi_master_sequencer    master_sequencer_D1308;
   svt_axi_master_sequencer    master_sequencer_D1309;
   svt_axi_master_sequencer    master_sequencer_D1310;
   svt_axi_master_sequencer    master_sequencer_D1311;
   svt_axi_master_sequencer    master_sequencer_D1312;
   svt_axi_master_sequencer    master_sequencer_D1313;
   svt_axi_master_sequencer    master_sequencer_D1314;
   svt_axi_master_sequencer    master_sequencer_D1315;
   svt_axi_master_sequencer    master_sequencer_D1316;
   svt_axi_master_sequencer    master_sequencer_D1317;
   svt_axi_master_sequencer    master_sequencer_D1318;
   svt_axi_master_sequencer    master_sequencer_D1319;
   svt_axi_master_sequencer    master_sequencer_D1320;
   svt_axi_master_sequencer    master_sequencer_D1321;
   svt_axi_master_sequencer    master_sequencer_D1322;
   svt_axi_master_sequencer    master_sequencer_D1323;
   svt_axi_master_sequencer    master_sequencer_D1324;
   svt_axi_master_sequencer    master_sequencer_D1325;
   svt_axi_master_sequencer    master_sequencer_D1326;
   svt_axi_master_sequencer    master_sequencer_D1327;
   svt_axi_master_sequencer    master_sequencer_D1328;
   svt_axi_master_sequencer    master_sequencer_D1329;
   svt_axi_master_sequencer    master_sequencer_D1330;
   svt_axi_master_sequencer    master_sequencer_D1331;
   svt_axi_master_sequencer    master_sequencer_D1332;
   svt_axi_master_sequencer    master_sequencer_D1333;
   svt_axi_master_sequencer    master_sequencer_D1334;
   svt_axi_master_sequencer    master_sequencer_D1335;
   svt_axi_master_sequencer    master_sequencer_D1336;
   svt_axi_master_sequencer    master_sequencer_D1337;
   svt_axi_master_sequencer    master_sequencer_D1338;
   svt_axi_master_sequencer    master_sequencer_D1339;
   svt_axi_master_sequencer    master_sequencer_D1340;
   svt_axi_master_sequencer    master_sequencer_D1341;
   svt_axi_master_sequencer    master_sequencer_D1342;
   svt_axi_master_sequencer    master_sequencer_D1343;
   svt_axi_master_sequencer    master_sequencer_D1344;
   svt_axi_master_sequencer    master_sequencer_D1345;
   svt_axi_master_sequencer    master_sequencer_D1346;
   svt_axi_master_sequencer    master_sequencer_D1347;
   svt_axi_master_sequencer    master_sequencer_D1348;
   svt_axi_master_sequencer    master_sequencer_D1349;
   svt_axi_master_sequencer    master_sequencer_D1350;
   svt_axi_master_sequencer    master_sequencer_D1351;
   svt_axi_master_sequencer    master_sequencer_D1352;
   svt_axi_master_sequencer    master_sequencer_D1353;
   svt_axi_master_sequencer    master_sequencer_D1354;
   svt_axi_master_sequencer    master_sequencer_D1355;
   svt_axi_master_sequencer    master_sequencer_D1356;
   svt_axi_master_sequencer    master_sequencer_D1357;
   svt_axi_master_sequencer    master_sequencer_D1358;
   svt_axi_master_sequencer    master_sequencer_D1359;
   svt_axi_master_sequencer    master_sequencer_D1360;
   svt_axi_master_sequencer    master_sequencer_D1361;
   svt_axi_master_sequencer    master_sequencer_D1362;
   svt_axi_master_sequencer    master_sequencer_D1363;
   svt_axi_master_sequencer    master_sequencer_D1364;
   svt_axi_master_sequencer    master_sequencer_D1365;
   svt_axi_master_sequencer    master_sequencer_D1366;
   svt_axi_master_sequencer    master_sequencer_D1367;
   svt_axi_master_sequencer    master_sequencer_D1368;
   svt_axi_master_sequencer    master_sequencer_D1369;
   svt_axi_master_sequencer    master_sequencer_D1370;
   svt_axi_master_sequencer    master_sequencer_D1371;
   svt_axi_master_sequencer    master_sequencer_D1372;
   svt_axi_master_sequencer    master_sequencer_D1373;
   svt_axi_master_sequencer    master_sequencer_D1374;
   svt_axi_master_sequencer    master_sequencer_D1375;
   svt_axi_master_sequencer    master_sequencer_D1376;
   svt_axi_master_sequencer    master_sequencer_D1377;
   svt_axi_master_sequencer    master_sequencer_D1378;
   svt_axi_master_sequencer    master_sequencer_D1379;
   svt_axi_master_sequencer    master_sequencer_D1380;
   svt_axi_master_sequencer    master_sequencer_D1381;
   svt_axi_master_sequencer    master_sequencer_D1382;
   svt_axi_master_sequencer    master_sequencer_D1383;
   svt_axi_master_sequencer    master_sequencer_D1384;
   svt_axi_master_sequencer    master_sequencer_D1385;
   svt_axi_master_sequencer    master_sequencer_D1386;
   svt_axi_master_sequencer    master_sequencer_D1387;
   svt_axi_master_sequencer    master_sequencer_D1388;
   svt_axi_master_sequencer    master_sequencer_D1389;
   svt_axi_master_sequencer    master_sequencer_D1390;
   svt_axi_master_sequencer    master_sequencer_D1391;
   svt_axi_master_sequencer    master_sequencer_D1392;
   svt_axi_master_sequencer    master_sequencer_D1393;
   svt_axi_master_sequencer    master_sequencer_D1394;
   svt_axi_master_sequencer    master_sequencer_D1395;
   svt_axi_master_sequencer    master_sequencer_D1396;
   svt_axi_master_sequencer    master_sequencer_D1397;
   svt_axi_master_sequencer    master_sequencer_D1398;
   svt_axi_master_sequencer    master_sequencer_D1399;
   svt_axi_master_sequencer    master_sequencer_D1400;
   svt_axi_master_sequencer    master_sequencer_D1401;
   svt_axi_master_sequencer    master_sequencer_D1402;
   svt_axi_master_sequencer    master_sequencer_D1403;
   svt_axi_master_sequencer    master_sequencer_D1404;
   svt_axi_master_sequencer    master_sequencer_D1405;
   svt_axi_master_sequencer    master_sequencer_D1406;
   svt_axi_master_sequencer    master_sequencer_D1407;
   svt_axi_master_sequencer    master_sequencer_D1408;
   svt_axi_master_sequencer    master_sequencer_D1409;
   svt_axi_master_sequencer    master_sequencer_D1410;
   svt_axi_master_sequencer    master_sequencer_D1411;
   svt_axi_master_sequencer    master_sequencer_D1412;
   svt_axi_master_sequencer    master_sequencer_D1413;
   svt_axi_master_sequencer    master_sequencer_D1414;
   svt_axi_master_sequencer    master_sequencer_D1415;
   svt_axi_master_sequencer    master_sequencer_D1416;
   svt_axi_master_sequencer    master_sequencer_D1417;
   svt_axi_master_sequencer    master_sequencer_D1418;
   svt_axi_master_sequencer    master_sequencer_D1419;
   svt_axi_master_sequencer    master_sequencer_D1420;
   svt_axi_master_sequencer    master_sequencer_D1421;
   svt_axi_master_sequencer    master_sequencer_D1422;
   svt_axi_master_sequencer    master_sequencer_D1423;
   svt_axi_master_sequencer    master_sequencer_D1424;
   svt_axi_master_sequencer    master_sequencer_D1425;
   svt_axi_master_sequencer    master_sequencer_D1426;
   svt_axi_master_sequencer    master_sequencer_D1427;
   svt_axi_master_sequencer    master_sequencer_D1428;
   svt_axi_master_sequencer    master_sequencer_D1429;
   svt_axi_master_sequencer    master_sequencer_D1430;
   svt_axi_master_sequencer    master_sequencer_D1431;
   svt_axi_master_sequencer    master_sequencer_D1432;
   svt_axi_master_sequencer    master_sequencer_D1433;
   svt_axi_master_sequencer    master_sequencer_D1434;
   svt_axi_master_sequencer    master_sequencer_D1435;
   svt_axi_master_sequencer    master_sequencer_D1436;
   svt_axi_master_sequencer    master_sequencer_D1437;
   svt_axi_master_sequencer    master_sequencer_D1438;
   svt_axi_master_sequencer    master_sequencer_D1439;
   svt_axi_master_sequencer    master_sequencer_D1440;
   svt_axi_master_sequencer    master_sequencer_D1441;
   svt_axi_master_sequencer    master_sequencer_D1442;
   svt_axi_master_sequencer    master_sequencer_D1443;
   svt_axi_master_sequencer    master_sequencer_D1444;
   svt_axi_master_sequencer    master_sequencer_D1445;
   svt_axi_master_sequencer    master_sequencer_D1446;
   svt_axi_master_sequencer    master_sequencer_D1447;
   svt_axi_master_sequencer    master_sequencer_D1448;
   svt_axi_master_sequencer    master_sequencer_D1449;
   svt_axi_master_sequencer    master_sequencer_D1450;
   svt_axi_master_sequencer    master_sequencer_D1451;
   svt_axi_master_sequencer    master_sequencer_D1452;
   svt_axi_master_sequencer    master_sequencer_D1453;
   svt_axi_master_sequencer    master_sequencer_D1454;
   svt_axi_master_sequencer    master_sequencer_D1455;
   svt_axi_master_sequencer    master_sequencer_D1456;
   svt_axi_master_sequencer    master_sequencer_D1457;
   svt_axi_master_sequencer    master_sequencer_D1458;
   svt_axi_master_sequencer    master_sequencer_D1459;
   svt_axi_master_sequencer    master_sequencer_D1460;
   svt_axi_master_sequencer    master_sequencer_D1461;
   svt_axi_master_sequencer    master_sequencer_D1462;
   svt_axi_master_sequencer    master_sequencer_D1463;
   svt_axi_master_sequencer    master_sequencer_D1464;
   svt_axi_master_sequencer    master_sequencer_D1465;
   svt_axi_master_sequencer    master_sequencer_D1466;
   svt_axi_master_sequencer    master_sequencer_D1467;
   svt_axi_master_sequencer    master_sequencer_D1468;
   svt_axi_master_sequencer    master_sequencer_D1469;
   svt_axi_master_sequencer    master_sequencer_D1470;
   svt_axi_master_sequencer    master_sequencer_D1471;
   svt_axi_master_sequencer    master_sequencer_D1472;
   svt_axi_master_sequencer    master_sequencer_D1473;
   svt_axi_master_sequencer    master_sequencer_D1474;
   svt_axi_master_sequencer    master_sequencer_D1475;
   svt_axi_master_sequencer    master_sequencer_D1476;
   svt_axi_master_sequencer    master_sequencer_D1477;
   svt_axi_master_sequencer    master_sequencer_D1478;
   svt_axi_master_sequencer    master_sequencer_D1479;
   svt_axi_master_sequencer    master_sequencer_D1480;
   svt_axi_master_sequencer    master_sequencer_D1481;
   svt_axi_master_sequencer    master_sequencer_D1482;
   svt_axi_master_sequencer    master_sequencer_D1483;
   svt_axi_master_sequencer    master_sequencer_D1484;
   svt_axi_master_sequencer    master_sequencer_D1485;
   svt_axi_master_sequencer    master_sequencer_D1486;
   svt_axi_master_sequencer    master_sequencer_D1487;
   svt_axi_master_sequencer    master_sequencer_D1488;
   svt_axi_master_sequencer    master_sequencer_D1489;
   svt_axi_master_sequencer    master_sequencer_D1490;
   svt_axi_master_sequencer    master_sequencer_D1491;
   svt_axi_master_sequencer    master_sequencer_D1492;
   svt_axi_master_sequencer    master_sequencer_D1493;
   svt_axi_master_sequencer    master_sequencer_D1494;
   svt_axi_master_sequencer    master_sequencer_D1495;
   svt_axi_master_sequencer    master_sequencer_D1496;
   svt_axi_master_sequencer    master_sequencer_D1497;
   svt_axi_master_sequencer    master_sequencer_D1498;
   svt_axi_master_sequencer    master_sequencer_D1499;
   svt_axi_master_sequencer    master_sequencer_D1500;
   svt_axi_master_sequencer    master_sequencer_D1501;
   svt_axi_master_sequencer    master_sequencer_D1502;
   svt_axi_master_sequencer    master_sequencer_D1503;
   svt_axi_master_sequencer    master_sequencer_D1504;
   svt_axi_master_sequencer    master_sequencer_D1505;
   svt_axi_master_sequencer    master_sequencer_D1506;
   svt_axi_master_sequencer    master_sequencer_D1507;
   svt_axi_master_sequencer    master_sequencer_D1508;
   svt_axi_master_sequencer    master_sequencer_D1509;
   svt_axi_master_sequencer    master_sequencer_D1510;
   svt_axi_master_sequencer    master_sequencer_D1511;
   svt_axi_master_sequencer    master_sequencer_D1512;
   svt_axi_master_sequencer    master_sequencer_D1513;
   svt_axi_master_sequencer    master_sequencer_D1514;
   svt_axi_master_sequencer    master_sequencer_D1515;
   svt_axi_master_sequencer    master_sequencer_D1516;
   svt_axi_master_sequencer    master_sequencer_D1517;
   svt_axi_master_sequencer    master_sequencer_D1518;
   svt_axi_master_sequencer    master_sequencer_D1519;
   svt_axi_master_sequencer    master_sequencer_D1520;
   svt_axi_master_sequencer    master_sequencer_D1521;
   svt_axi_master_sequencer    master_sequencer_D1522;
   svt_axi_master_sequencer    master_sequencer_D1523;
   svt_axi_master_sequencer    master_sequencer_D1524;
   svt_axi_master_sequencer    master_sequencer_D1525;
   svt_axi_master_sequencer    master_sequencer_D1526;
   svt_axi_master_sequencer    master_sequencer_D1527;
   svt_axi_master_sequencer    master_sequencer_D1528;
   svt_axi_master_sequencer    master_sequencer_D1529;
   svt_axi_master_sequencer    master_sequencer_D1530;
   svt_axi_master_sequencer    master_sequencer_D1531;
   svt_axi_master_sequencer    master_sequencer_D1532;
   svt_axi_master_sequencer    master_sequencer_D1533;
   svt_axi_master_sequencer    master_sequencer_D1534;
   svt_axi_master_sequencer    master_sequencer_D1535;
   svt_axi_master_sequencer    master_sequencer_D1536;
   svt_axi_master_sequencer    master_sequencer_D1537;
   svt_axi_master_sequencer    master_sequencer_D1538;
   svt_axi_master_sequencer    master_sequencer_D1539;
   svt_axi_master_sequencer    master_sequencer_D1540;
   svt_axi_master_sequencer    master_sequencer_D1541;
   svt_axi_master_sequencer    master_sequencer_D1542;
   svt_axi_master_sequencer    master_sequencer_D1543;
   svt_axi_master_sequencer    master_sequencer_D1544;
   svt_axi_master_sequencer    master_sequencer_D1545;
   svt_axi_master_sequencer    master_sequencer_D1546;
   svt_axi_master_sequencer    master_sequencer_D1547;
   svt_axi_master_sequencer    master_sequencer_D1548;
   svt_axi_master_sequencer    master_sequencer_D1549;
   svt_axi_master_sequencer    master_sequencer_D1550;
   svt_axi_master_sequencer    master_sequencer_D1551;
   svt_axi_master_sequencer    master_sequencer_D1552;
   svt_axi_master_sequencer    master_sequencer_D1553;
   svt_axi_master_sequencer    master_sequencer_D1554;
   svt_axi_master_sequencer    master_sequencer_D1555;
   svt_axi_master_sequencer    master_sequencer_D1556;
   svt_axi_master_sequencer    master_sequencer_D1557;
   svt_axi_master_sequencer    master_sequencer_D1558;
   svt_axi_master_sequencer    master_sequencer_D1559;
   svt_axi_master_sequencer    master_sequencer_D1560;
   svt_axi_master_sequencer    master_sequencer_D1561;
   svt_axi_master_sequencer    master_sequencer_D1562;
   svt_axi_master_sequencer    master_sequencer_D1563;
   svt_axi_master_sequencer    master_sequencer_D1564;
   svt_axi_master_sequencer    master_sequencer_D1565;
   svt_axi_master_sequencer    master_sequencer_D1566;
   svt_axi_master_sequencer    master_sequencer_D1567;
   svt_axi_master_sequencer    master_sequencer_D1568;
   svt_axi_master_sequencer    master_sequencer_D1569;
   svt_axi_master_sequencer    master_sequencer_D1570;
   svt_axi_master_sequencer    master_sequencer_D1571;
   svt_axi_master_sequencer    master_sequencer_D1572;
   svt_axi_master_sequencer    master_sequencer_D1573;
   svt_axi_master_sequencer    master_sequencer_D1574;
   svt_axi_master_sequencer    master_sequencer_D1575;
   svt_axi_master_sequencer    master_sequencer_D1576;
   svt_axi_master_sequencer    master_sequencer_D1577;
   svt_axi_master_sequencer    master_sequencer_D1578;
   svt_axi_master_sequencer    master_sequencer_D1579;
   svt_axi_master_sequencer    master_sequencer_D1580;
   svt_axi_master_sequencer    master_sequencer_D1581;
   svt_axi_master_sequencer    master_sequencer_D1582;
   svt_axi_master_sequencer    master_sequencer_D1583;
   svt_axi_master_sequencer    master_sequencer_D1584;
   svt_axi_master_sequencer    master_sequencer_D1585;
   svt_axi_master_sequencer    master_sequencer_D1586;
   svt_axi_master_sequencer    master_sequencer_D1587;
   svt_axi_master_sequencer    master_sequencer_D1588;
   svt_axi_master_sequencer    master_sequencer_D1589;
   svt_axi_master_sequencer    master_sequencer_D1590;
   svt_axi_master_sequencer    master_sequencer_D1591;
   svt_axi_master_sequencer    master_sequencer_D1592;
   svt_axi_master_sequencer    master_sequencer_D1593;
   svt_axi_master_sequencer    master_sequencer_D1594;
   svt_axi_master_sequencer    master_sequencer_D1595;
   svt_axi_master_sequencer    master_sequencer_D1596;
   svt_axi_master_sequencer    master_sequencer_D1597;
   svt_axi_master_sequencer    master_sequencer_D1598;
   svt_axi_master_sequencer    master_sequencer_D1599;
   svt_axi_master_sequencer    master_sequencer_D1600;
   svt_axi_master_sequencer    master_sequencer_D1601;
   svt_axi_master_sequencer    master_sequencer_D1602;
   svt_axi_master_sequencer    master_sequencer_D1603;
   svt_axi_master_sequencer    master_sequencer_D1604;
   svt_axi_master_sequencer    master_sequencer_D1605;
   svt_axi_master_sequencer    master_sequencer_D1606;
   svt_axi_master_sequencer    master_sequencer_D1607;
   svt_axi_master_sequencer    master_sequencer_D1608;
   svt_axi_master_sequencer    master_sequencer_D1609;
   svt_axi_master_sequencer    master_sequencer_D1610;
   svt_axi_master_sequencer    master_sequencer_D1611;
   svt_axi_master_sequencer    master_sequencer_D1612;
   svt_axi_master_sequencer    master_sequencer_D1613;
   svt_axi_master_sequencer    master_sequencer_D1614;
   svt_axi_master_sequencer    master_sequencer_D1615;
   svt_axi_master_sequencer    master_sequencer_D1616;
   svt_axi_master_sequencer    master_sequencer_D1617;
   svt_axi_master_sequencer    master_sequencer_D1618;
   svt_axi_master_sequencer    master_sequencer_D1619;
   svt_axi_master_sequencer    master_sequencer_D1620;
   svt_axi_master_sequencer    master_sequencer_D1621;
   svt_axi_master_sequencer    master_sequencer_D1622;
   svt_axi_master_sequencer    master_sequencer_D1623;
   svt_axi_master_sequencer    master_sequencer_D1624;
   svt_axi_master_sequencer    master_sequencer_D1625;
   svt_axi_master_sequencer    master_sequencer_D1626;
   svt_axi_master_sequencer    master_sequencer_D1627;
   svt_axi_master_sequencer    master_sequencer_D1628;
   svt_axi_master_sequencer    master_sequencer_D1629;
   svt_axi_master_sequencer    master_sequencer_D1630;
   svt_axi_master_sequencer    master_sequencer_D1631;
   svt_axi_master_sequencer    master_sequencer_D1632;
   svt_axi_master_sequencer    master_sequencer_D1633;
   svt_axi_master_sequencer    master_sequencer_D1634;
   svt_axi_master_sequencer    master_sequencer_D1635;
   svt_axi_master_sequencer    master_sequencer_D1636;
   svt_axi_master_sequencer    master_sequencer_D1637;
   svt_axi_master_sequencer    master_sequencer_D1638;
   svt_axi_master_sequencer    master_sequencer_D1639;
   svt_axi_master_sequencer    master_sequencer_D1640;
   svt_axi_master_sequencer    master_sequencer_D1641;
   svt_axi_master_sequencer    master_sequencer_D1642;
   svt_axi_master_sequencer    master_sequencer_D1643;
   svt_axi_master_sequencer    master_sequencer_D1644;
   svt_axi_master_sequencer    master_sequencer_D1645;
   svt_axi_master_sequencer    master_sequencer_D1646;
   svt_axi_master_sequencer    master_sequencer_D1647;
   svt_axi_master_sequencer    master_sequencer_D1648;
   svt_axi_master_sequencer    master_sequencer_D1649;
   svt_axi_master_sequencer    master_sequencer_D1650;
   svt_axi_master_sequencer    master_sequencer_D1651;
   svt_axi_master_sequencer    master_sequencer_D1652;
   svt_axi_master_sequencer    master_sequencer_D1653;
   svt_axi_master_sequencer    master_sequencer_D1654;
   svt_axi_master_sequencer    master_sequencer_D1655;
   svt_axi_master_sequencer    master_sequencer_D1656;
   svt_axi_master_sequencer    master_sequencer_D1657;
   svt_axi_master_sequencer    master_sequencer_D1658;
   svt_axi_master_sequencer    master_sequencer_D1659;
   svt_axi_master_sequencer    master_sequencer_D1660;
   svt_axi_master_sequencer    master_sequencer_D1661;
   svt_axi_master_sequencer    master_sequencer_D1662;
   svt_axi_master_sequencer    master_sequencer_D1663;
   svt_axi_master_sequencer    master_sequencer_D1664;
   svt_axi_master_sequencer    master_sequencer_D1665;
   svt_axi_master_sequencer    master_sequencer_D1666;
   svt_axi_master_sequencer    master_sequencer_D1667;
   svt_axi_master_sequencer    master_sequencer_D1668;
   svt_axi_master_sequencer    master_sequencer_D1669;
   svt_axi_master_sequencer    master_sequencer_D1670;
   svt_axi_master_sequencer    master_sequencer_D1671;
   svt_axi_master_sequencer    master_sequencer_D1672;
   svt_axi_master_sequencer    master_sequencer_D1673;
   svt_axi_master_sequencer    master_sequencer_D1674;
   svt_axi_master_sequencer    master_sequencer_D1675;
   svt_axi_master_sequencer    master_sequencer_D1676;
   svt_axi_master_sequencer    master_sequencer_D1677;
   svt_axi_master_sequencer    master_sequencer_D1678;
   svt_axi_master_sequencer    master_sequencer_D1679;
   svt_axi_master_sequencer    master_sequencer_D1680;
   svt_axi_master_sequencer    master_sequencer_D1681;
   svt_axi_master_sequencer    master_sequencer_D1682;
   svt_axi_master_sequencer    master_sequencer_D1683;
   svt_axi_master_sequencer    master_sequencer_D1684;
   svt_axi_master_sequencer    master_sequencer_D1685;
   svt_axi_master_sequencer    master_sequencer_D1686;
   svt_axi_master_sequencer    master_sequencer_D1687;
   svt_axi_master_sequencer    master_sequencer_D1688;
   svt_axi_master_sequencer    master_sequencer_D1689;
   svt_axi_master_sequencer    master_sequencer_D1690;
   svt_axi_master_sequencer    master_sequencer_D1691;
   svt_axi_master_sequencer    master_sequencer_D1692;
   svt_axi_master_sequencer    master_sequencer_D1693;
   svt_axi_master_sequencer    master_sequencer_D1694;
   svt_axi_master_sequencer    master_sequencer_D1695;
   svt_axi_master_sequencer    master_sequencer_D1696;
   svt_axi_master_sequencer    master_sequencer_D1697;
   svt_axi_master_sequencer    master_sequencer_D1698;
   svt_axi_master_sequencer    master_sequencer_D1699;
   svt_axi_master_sequencer    master_sequencer_D1700;
   svt_axi_master_sequencer    master_sequencer_D1701;
   svt_axi_master_sequencer    master_sequencer_D1702;
   svt_axi_master_sequencer    master_sequencer_D1703;
   svt_axi_master_sequencer    master_sequencer_D1704;
   svt_axi_master_sequencer    master_sequencer_D1705;
   svt_axi_master_sequencer    master_sequencer_D1706;
   svt_axi_master_sequencer    master_sequencer_D1707;
   svt_axi_master_sequencer    master_sequencer_D1708;
   svt_axi_master_sequencer    master_sequencer_D1709;
   svt_axi_master_sequencer    master_sequencer_D1710;
   svt_axi_master_sequencer    master_sequencer_D1711;
   svt_axi_master_sequencer    master_sequencer_D1712;
   svt_axi_master_sequencer    master_sequencer_D1713;
   svt_axi_master_sequencer    master_sequencer_D1714;
   svt_axi_master_sequencer    master_sequencer_D1715;
   svt_axi_master_sequencer    master_sequencer_D1716;
   svt_axi_master_sequencer    master_sequencer_D1717;
   svt_axi_master_sequencer    master_sequencer_D1718;
   svt_axi_master_sequencer    master_sequencer_D1719;
   svt_axi_master_sequencer    master_sequencer_D1720;
   svt_axi_master_sequencer    master_sequencer_D1721;
   svt_axi_master_sequencer    master_sequencer_D1722;
   svt_axi_master_sequencer    master_sequencer_D1723;
   svt_axi_master_sequencer    master_sequencer_D1724;
   svt_axi_master_sequencer    master_sequencer_D1725;
   svt_axi_master_sequencer    master_sequencer_D1726;
   svt_axi_master_sequencer    master_sequencer_D1727;
   svt_axi_master_sequencer    master_sequencer_D1728;
   svt_axi_master_sequencer    master_sequencer_D1729;
   svt_axi_master_sequencer    master_sequencer_D1730;
   svt_axi_master_sequencer    master_sequencer_D1731;
   svt_axi_master_sequencer    master_sequencer_D1732;
   svt_axi_master_sequencer    master_sequencer_D1733;
   svt_axi_master_sequencer    master_sequencer_D1734;
   svt_axi_master_sequencer    master_sequencer_D1735;
   svt_axi_master_sequencer    master_sequencer_D1736;
   svt_axi_master_sequencer    master_sequencer_D1737;
   svt_axi_master_sequencer    master_sequencer_D1738;
   svt_axi_master_sequencer    master_sequencer_D1739;
   svt_axi_master_sequencer    master_sequencer_D1740;
   svt_axi_master_sequencer    master_sequencer_D1741;
   svt_axi_master_sequencer    master_sequencer_D1742;
   svt_axi_master_sequencer    master_sequencer_D1743;
   svt_axi_master_sequencer    master_sequencer_D1744;
   svt_axi_master_sequencer    master_sequencer_D1745;
   svt_axi_master_sequencer    master_sequencer_D1746;
   svt_axi_master_sequencer    master_sequencer_D1747;
   svt_axi_master_sequencer    master_sequencer_D1748;
   svt_axi_master_sequencer    master_sequencer_D1749;
   svt_axi_master_sequencer    master_sequencer_D1750;
   svt_axi_master_sequencer    master_sequencer_D1751;
   svt_axi_master_sequencer    master_sequencer_D1752;
   svt_axi_master_sequencer    master_sequencer_D1753;
   svt_axi_master_sequencer    master_sequencer_D1754;
   svt_axi_master_sequencer    master_sequencer_D1755;
   svt_axi_master_sequencer    master_sequencer_D1756;
   svt_axi_master_sequencer    master_sequencer_D1757;
   svt_axi_master_sequencer    master_sequencer_D1758;
   svt_axi_master_sequencer    master_sequencer_D1759;
   svt_axi_master_sequencer    master_sequencer_D1760;
   svt_axi_master_sequencer    master_sequencer_D1761;
   svt_axi_master_sequencer    master_sequencer_D1762;
   svt_axi_master_sequencer    master_sequencer_D1763;
   svt_axi_master_sequencer    master_sequencer_D1764;
   svt_axi_master_sequencer    master_sequencer_D1765;
   svt_axi_master_sequencer    master_sequencer_D1766;
   svt_axi_master_sequencer    master_sequencer_D1767;
   svt_axi_master_sequencer    master_sequencer_D1768;
   svt_axi_master_sequencer    master_sequencer_D1769;
   svt_axi_master_sequencer    master_sequencer_D1770;
   svt_axi_master_sequencer    master_sequencer_D1771;
   svt_axi_master_sequencer    master_sequencer_D1772;
   svt_axi_master_sequencer    master_sequencer_D1773;
   svt_axi_master_sequencer    master_sequencer_D1774;
   svt_axi_master_sequencer    master_sequencer_D1775;
   svt_axi_master_sequencer    master_sequencer_D1776;
   svt_axi_master_sequencer    master_sequencer_D1777;
   svt_axi_master_sequencer    master_sequencer_D1778;
   svt_axi_master_sequencer    master_sequencer_D1779;
   svt_axi_master_sequencer    master_sequencer_D1780;
   svt_axi_master_sequencer    master_sequencer_D1781;
   svt_axi_master_sequencer    master_sequencer_D1782;
   svt_axi_master_sequencer    master_sequencer_D1783;
   svt_axi_master_sequencer    master_sequencer_D1784;
   svt_axi_master_sequencer    master_sequencer_D1785;
   svt_axi_master_sequencer    master_sequencer_D1786;
   svt_axi_master_sequencer    master_sequencer_D1787;
   svt_axi_master_sequencer    master_sequencer_D1788;
   svt_axi_master_sequencer    master_sequencer_D1789;
   svt_axi_master_sequencer    master_sequencer_D1790;
   svt_axi_master_sequencer    master_sequencer_D1791;
   svt_axi_master_sequencer    master_sequencer_D1792;
   svt_axi_master_sequencer    master_sequencer_D1793;
   svt_axi_master_sequencer    master_sequencer_D1794;
   svt_axi_master_sequencer    master_sequencer_D1795;
   svt_axi_master_sequencer    master_sequencer_D1796;
   svt_axi_master_sequencer    master_sequencer_D1797;
   svt_axi_master_sequencer    master_sequencer_D1798;
   svt_axi_master_sequencer    master_sequencer_D1799;
   svt_axi_master_sequencer    master_sequencer_D1800;
   svt_axi_master_sequencer    master_sequencer_D1801;
   svt_axi_master_sequencer    master_sequencer_D1802;
   svt_axi_master_sequencer    master_sequencer_D1803;
   svt_axi_master_sequencer    master_sequencer_D1804;
   svt_axi_master_sequencer    master_sequencer_D1805;
   svt_axi_master_sequencer    master_sequencer_D1806;
   svt_axi_master_sequencer    master_sequencer_D1807;
   svt_axi_master_sequencer    master_sequencer_D1808;
   svt_axi_master_sequencer    master_sequencer_D1809;
   svt_axi_master_sequencer    master_sequencer_D1810;
   svt_axi_master_sequencer    master_sequencer_D1811;
   svt_axi_master_sequencer    master_sequencer_D1812;
   svt_axi_master_sequencer    master_sequencer_D1813;
   svt_axi_master_sequencer    master_sequencer_D1814;
   svt_axi_master_sequencer    master_sequencer_D1815;
   svt_axi_master_sequencer    master_sequencer_D1816;
   svt_axi_master_sequencer    master_sequencer_D1817;
   svt_axi_master_sequencer    master_sequencer_D1818;
   svt_axi_master_sequencer    master_sequencer_D1819;
   svt_axi_master_sequencer    master_sequencer_D1820;
   svt_axi_master_sequencer    master_sequencer_D1821;
   svt_axi_master_sequencer    master_sequencer_D1822;
   svt_axi_master_sequencer    master_sequencer_D1823;
   svt_axi_master_sequencer    master_sequencer_D1824;
   svt_axi_master_sequencer    master_sequencer_D1825;
   svt_axi_master_sequencer    master_sequencer_D1826;
   svt_axi_master_sequencer    master_sequencer_D1827;
   svt_axi_master_sequencer    master_sequencer_D1828;
   svt_axi_master_sequencer    master_sequencer_D1829;
   svt_axi_master_sequencer    master_sequencer_D1830;
   svt_axi_master_sequencer    master_sequencer_D1831;
   svt_axi_master_sequencer    master_sequencer_D1832;
   svt_axi_master_sequencer    master_sequencer_D1833;
   svt_axi_master_sequencer    master_sequencer_D1834;
   svt_axi_master_sequencer    master_sequencer_D1835;
   svt_axi_master_sequencer    master_sequencer_D1836;
   svt_axi_master_sequencer    master_sequencer_D1837;
   svt_axi_master_sequencer    master_sequencer_D1838;
   svt_axi_master_sequencer    master_sequencer_D1839;
   svt_axi_master_sequencer    master_sequencer_D1840;
   svt_axi_master_sequencer    master_sequencer_D1841;
   svt_axi_master_sequencer    master_sequencer_D1842;
   svt_axi_master_sequencer    master_sequencer_D1843;
   svt_axi_master_sequencer    master_sequencer_D1844;
   svt_axi_master_sequencer    master_sequencer_D1845;
   svt_axi_master_sequencer    master_sequencer_D1846;
   svt_axi_master_sequencer    master_sequencer_D1847;
   svt_axi_master_sequencer    master_sequencer_D1848;
   svt_axi_master_sequencer    master_sequencer_D1849;
   svt_axi_master_sequencer    master_sequencer_D1850;
   svt_axi_master_sequencer    master_sequencer_D1851;
   svt_axi_master_sequencer    master_sequencer_D1852;
   svt_axi_master_sequencer    master_sequencer_D1853;
   svt_axi_master_sequencer    master_sequencer_D1854;
   svt_axi_master_sequencer    master_sequencer_D1855;
   svt_axi_master_sequencer    master_sequencer_D1856;
   svt_axi_master_sequencer    master_sequencer_D1857;
   svt_axi_master_sequencer    master_sequencer_D1858;
   svt_axi_master_sequencer    master_sequencer_D1859;
   svt_axi_master_sequencer    master_sequencer_D1860;
   svt_axi_master_sequencer    master_sequencer_D1861;
   svt_axi_master_sequencer    master_sequencer_D1862;
   svt_axi_master_sequencer    master_sequencer_D1863;
   svt_axi_master_sequencer    master_sequencer_D1864;
   svt_axi_master_sequencer    master_sequencer_D1865;
   svt_axi_master_sequencer    master_sequencer_D1866;
   svt_axi_master_sequencer    master_sequencer_D1867;
   svt_axi_master_sequencer    master_sequencer_D1868;
   svt_axi_master_sequencer    master_sequencer_D1869;
   svt_axi_master_sequencer    master_sequencer_D1870;
   svt_axi_master_sequencer    master_sequencer_D1871;
   svt_axi_master_sequencer    master_sequencer_D1872;
   svt_axi_master_sequencer    master_sequencer_D1873;
   svt_axi_master_sequencer    master_sequencer_D1874;
   svt_axi_master_sequencer    master_sequencer_D1875;
   svt_axi_master_sequencer    master_sequencer_D1876;
   svt_axi_master_sequencer    master_sequencer_D1877;
   svt_axi_master_sequencer    master_sequencer_D1878;
   svt_axi_master_sequencer    master_sequencer_D1879;
   svt_axi_master_sequencer    master_sequencer_D1880;
   svt_axi_master_sequencer    master_sequencer_D1881;
   svt_axi_master_sequencer    master_sequencer_D1882;
   svt_axi_master_sequencer    master_sequencer_D1883;
   svt_axi_master_sequencer    master_sequencer_D1884;
   svt_axi_master_sequencer    master_sequencer_D1885;
   svt_axi_master_sequencer    master_sequencer_D1886;
   svt_axi_master_sequencer    master_sequencer_D1887;
   svt_axi_master_sequencer    master_sequencer_D1888;
   svt_axi_master_sequencer    master_sequencer_D1889;
   svt_axi_master_sequencer    master_sequencer_D1890;
   svt_axi_master_sequencer    master_sequencer_D1891;
   svt_axi_master_sequencer    master_sequencer_D1892;
   svt_axi_master_sequencer    master_sequencer_D1893;
   svt_axi_master_sequencer    master_sequencer_D1894;
   svt_axi_master_sequencer    master_sequencer_D1895;
   svt_axi_master_sequencer    master_sequencer_D1896;
   svt_axi_master_sequencer    master_sequencer_D1897;
   svt_axi_master_sequencer    master_sequencer_D1898;
   svt_axi_master_sequencer    master_sequencer_D1899;
   svt_axi_master_sequencer    master_sequencer_D1900;
   svt_axi_master_sequencer    master_sequencer_D1901;
   svt_axi_master_sequencer    master_sequencer_D1902;
   svt_axi_master_sequencer    master_sequencer_D1903;
   svt_axi_master_sequencer    master_sequencer_D1904;
   svt_axi_master_sequencer    master_sequencer_D1905;
   svt_axi_master_sequencer    master_sequencer_D1906;
   svt_axi_master_sequencer    master_sequencer_D1907;
   svt_axi_master_sequencer    master_sequencer_D1908;
   svt_axi_master_sequencer    master_sequencer_D1909;
   svt_axi_master_sequencer    master_sequencer_D1910;
   svt_axi_master_sequencer    master_sequencer_D1911;
   svt_axi_master_sequencer    master_sequencer_D1912;
   svt_axi_master_sequencer    master_sequencer_D1913;
   svt_axi_master_sequencer    master_sequencer_D1914;
   svt_axi_master_sequencer    master_sequencer_D1915;
   svt_axi_master_sequencer    master_sequencer_D1916;
   svt_axi_master_sequencer    master_sequencer_D1917;
   svt_axi_master_sequencer    master_sequencer_D1918;
   svt_axi_master_sequencer    master_sequencer_D1919;
   svt_axi_master_sequencer    master_sequencer_D1920;
   svt_axi_master_sequencer    master_sequencer_D1921;
   svt_axi_master_sequencer    master_sequencer_D1922;
   svt_axi_master_sequencer    master_sequencer_D1923;
   svt_axi_master_sequencer    master_sequencer_D1924;
   svt_axi_master_sequencer    master_sequencer_D1925;
   svt_axi_master_sequencer    master_sequencer_D1926;
   svt_axi_master_sequencer    master_sequencer_D1927;
   svt_axi_master_sequencer    master_sequencer_D1928;
   svt_axi_master_sequencer    master_sequencer_D1929;
   svt_axi_master_sequencer    master_sequencer_D1930;
   svt_axi_master_sequencer    master_sequencer_D1931;
   svt_axi_master_sequencer    master_sequencer_D1932;
   svt_axi_master_sequencer    master_sequencer_D1933;
   svt_axi_master_sequencer    master_sequencer_D1934;
   svt_axi_master_sequencer    master_sequencer_D1935;
   svt_axi_master_sequencer    master_sequencer_D1936;
   svt_axi_master_sequencer    master_sequencer_D1937;
   svt_axi_master_sequencer    master_sequencer_D1938;
   svt_axi_master_sequencer    master_sequencer_D1939;
   svt_axi_master_sequencer    master_sequencer_D1940;
   svt_axi_master_sequencer    master_sequencer_D1941;
   svt_axi_master_sequencer    master_sequencer_D1942;
   svt_axi_master_sequencer    master_sequencer_D1943;
   svt_axi_master_sequencer    master_sequencer_D1944;
   svt_axi_master_sequencer    master_sequencer_D1945;
   svt_axi_master_sequencer    master_sequencer_D1946;
   svt_axi_master_sequencer    master_sequencer_D1947;
   svt_axi_master_sequencer    master_sequencer_D1948;
   svt_axi_master_sequencer    master_sequencer_D1949;
   svt_axi_master_sequencer    master_sequencer_D1950;
   svt_axi_master_sequencer    master_sequencer_D1951;
   svt_axi_master_sequencer    master_sequencer_D1952;
   svt_axi_master_sequencer    master_sequencer_D1953;
   svt_axi_master_sequencer    master_sequencer_D1954;
   svt_axi_master_sequencer    master_sequencer_D1955;
   svt_axi_master_sequencer    master_sequencer_D1956;
   svt_axi_master_sequencer    master_sequencer_D1957;
   svt_axi_master_sequencer    master_sequencer_D1958;
   svt_axi_master_sequencer    master_sequencer_D1959;
   svt_axi_master_sequencer    master_sequencer_D1960;
   svt_axi_master_sequencer    master_sequencer_D1961;
   svt_axi_master_sequencer    master_sequencer_D1962;
   svt_axi_master_sequencer    master_sequencer_D1963;
   svt_axi_master_sequencer    master_sequencer_D1964;
   svt_axi_master_sequencer    master_sequencer_D1965;
   svt_axi_master_sequencer    master_sequencer_D1966;
   svt_axi_master_sequencer    master_sequencer_D1967;
   svt_axi_master_sequencer    master_sequencer_D1968;
   svt_axi_master_sequencer    master_sequencer_D1969;
   svt_axi_master_sequencer    master_sequencer_D1970;
   svt_axi_master_sequencer    master_sequencer_D1971;
   svt_axi_master_sequencer    master_sequencer_D1972;
   svt_axi_master_sequencer    master_sequencer_D1973;
   svt_axi_master_sequencer    master_sequencer_D1974;
   svt_axi_master_sequencer    master_sequencer_D1975;
   svt_axi_master_sequencer    master_sequencer_D1976;
   svt_axi_master_sequencer    master_sequencer_D1977;
   svt_axi_master_sequencer    master_sequencer_D1978;
   svt_axi_master_sequencer    master_sequencer_D1979;
   svt_axi_master_sequencer    master_sequencer_D1980;
   svt_axi_master_sequencer    master_sequencer_D1981;
   svt_axi_master_sequencer    master_sequencer_D1982;
   svt_axi_master_sequencer    master_sequencer_D1983;
   svt_axi_master_sequencer    master_sequencer_D1984;
   svt_axi_master_sequencer    master_sequencer_D1985;
   svt_axi_master_sequencer    master_sequencer_D1986;
   svt_axi_master_sequencer    master_sequencer_D1987;
   svt_axi_master_sequencer    master_sequencer_D1988;
   svt_axi_master_sequencer    master_sequencer_D1989;
   svt_axi_master_sequencer    master_sequencer_D1990;
   svt_axi_master_sequencer    master_sequencer_D1991;
   svt_axi_master_sequencer    master_sequencer_D1992;
   svt_axi_master_sequencer    master_sequencer_D1993;
   svt_axi_master_sequencer    master_sequencer_D1994;
   svt_axi_master_sequencer    master_sequencer_D1995;
   svt_axi_master_sequencer    master_sequencer_D1996;
   svt_axi_master_sequencer    master_sequencer_D1997;
   svt_axi_master_sequencer    master_sequencer_D1998;
   svt_axi_master_sequencer    master_sequencer_D1999;
   svt_axi_master_sequencer    master_sequencer_D2000;
   svt_axi_master_sequencer    master_sequencer_D2001;
   svt_axi_master_sequencer    master_sequencer_D2002;
   svt_axi_master_sequencer    master_sequencer_D2003;
   svt_axi_master_sequencer    master_sequencer_D2004;
   svt_axi_master_sequencer    master_sequencer_D2005;
   svt_axi_master_sequencer    master_sequencer_D2006;
   svt_axi_master_sequencer    master_sequencer_D2007;
   svt_axi_master_sequencer    master_sequencer_D2008;
   svt_axi_master_sequencer    master_sequencer_D2009;
   svt_axi_master_sequencer    master_sequencer_D2010;
   svt_axi_master_sequencer    master_sequencer_D2011;
   svt_axi_master_sequencer    master_sequencer_D2012;
   svt_axi_master_sequencer    master_sequencer_D2013;
   svt_axi_master_sequencer    master_sequencer_D2014;
   svt_axi_master_sequencer    master_sequencer_D2015;
   svt_axi_master_sequencer    master_sequencer_D2016;
   svt_axi_master_sequencer    master_sequencer_D2017;
   svt_axi_master_sequencer    master_sequencer_D2018;
   svt_axi_master_sequencer    master_sequencer_D2019;
   svt_axi_master_sequencer    master_sequencer_D2020;
   svt_axi_master_sequencer    master_sequencer_D2021;
   svt_axi_master_sequencer    master_sequencer_D2022;
   svt_axi_master_sequencer    master_sequencer_D2023;
   svt_axi_master_sequencer    master_sequencer_D2024;
   svt_axi_master_sequencer    master_sequencer_D2025;
   svt_axi_master_sequencer    master_sequencer_D2026;
   svt_axi_master_sequencer    master_sequencer_D2027;
   svt_axi_master_sequencer    master_sequencer_D2028;
   svt_axi_master_sequencer    master_sequencer_D2029;
   svt_axi_master_sequencer    master_sequencer_D2030;
   svt_axi_master_sequencer    master_sequencer_D2031;
   svt_axi_master_sequencer    master_sequencer_D2032;
   svt_axi_master_sequencer    master_sequencer_D2033;
   svt_axi_master_sequencer    master_sequencer_D2034;
   svt_axi_master_sequencer    master_sequencer_D2035;
   svt_axi_master_sequencer    master_sequencer_D2036;
   svt_axi_master_sequencer    master_sequencer_D2037;
   svt_axi_master_sequencer    master_sequencer_D2038;
   svt_axi_master_sequencer    master_sequencer_D2039;
   svt_axi_master_sequencer    master_sequencer_D2040;
   svt_axi_master_sequencer    master_sequencer_D2041;
   svt_axi_master_sequencer    master_sequencer_D2042;
   svt_axi_master_sequencer    master_sequencer_D2043;
   svt_axi_master_sequencer    master_sequencer_D2044;
   svt_axi_master_sequencer    master_sequencer_D2045;
   svt_axi_master_sequencer    master_sequencer_D2046;
   svt_axi_master_sequencer    master_sequencer_D2047;
   `endif


  function new(string name="pf_vf_mux_virtual_sequencer", uvm_component parent=null);
    super.new(name,parent);
  endfunction // new


  virtual function void build_phase(uvm_phase phase);
    `uvm_info("build_phase", "Entered...", UVM_LOW)

    super.build_phase(phase);

    if (!uvm_config_db#(AXI_RESET_MP)::get(this, "", "reset_mp", reset_mp)) begin
      `uvm_fatal("build_phase", "An axi_reset_modport must be set using the config db.");
    end

    `uvm_info("build_phase", "Exiting...", UVM_LOW)
  endfunction

endclass

`endif // GUARD_pf_vf_mux_virtual_sequencer_SV
