// Copyright (C) 2020 Intel Corporation
// SPDX-License-Identifier: MIT

// avst_pipeline_st_pipeline_stage_0.v

// Generated using ACDS version 22.1 174

`timescale 1 ps / 1 ps
module avst_pipeline_st_pipeline_stage_0 #(
		parameter SYMBOLS_PER_BEAT = 64,
		parameter BITS_PER_SYMBOL  = 8,
		parameter USE_PACKETS      = 1,
		parameter USE_EMPTY        = 1,
		parameter EMPTY_WIDTH      = 6,
		parameter CHANNEL_WIDTH    = 0,
		parameter PACKET_WIDTH     = 2,
		parameter ERROR_WIDTH      = 1,
		parameter PIPELINE_READY   = 1,
		parameter SYNC_RESET       = 1
	) (
		input  wire         clk,               //       cr0.clk
		input  wire         reset,             // cr0_reset.reset
		output wire         in_ready,          //     sink0.ready
		input  wire         in_valid,          //          .valid
		input  wire         in_startofpacket,  //          .startofpacket
		input  wire         in_endofpacket,    //          .endofpacket
		input  wire [5:0]   in_empty,          //          .empty
		input  wire [0:0]   in_error,          //          .error
		input  wire [511:0] in_data,           //          .data
		input  wire         out_ready,         //   source0.ready
		output wire         out_valid,         //          .valid
		output wire         out_startofpacket, //          .startofpacket
		output wire         out_endofpacket,   //          .endofpacket
		output wire [5:0]   out_empty,         //          .empty
		output wire [0:0]   out_error,         //          .error
		output wire [511:0] out_data           //          .data
	);

	avst_pipeline_st_pipeline_stage_0_altera_avalon_st_pipeline_stage_1920_zterisq #(
		.SYMBOLS_PER_BEAT (SYMBOLS_PER_BEAT),
		.BITS_PER_SYMBOL  (BITS_PER_SYMBOL),
		.USE_PACKETS      (USE_PACKETS),
		.USE_EMPTY        (USE_EMPTY),
		.EMPTY_WIDTH      (EMPTY_WIDTH),
		.CHANNEL_WIDTH    (CHANNEL_WIDTH),
		.PACKET_WIDTH     (PACKET_WIDTH),
		.ERROR_WIDTH      (ERROR_WIDTH),
		.PIPELINE_READY   (PIPELINE_READY),
		.SYNC_RESET       (SYNC_RESET)
	) st_pipeline_stage_0 (
		.clk               (clk),               //   input,    width = 1,       cr0.clk
		.reset             (reset),             //   input,    width = 1, cr0_reset.reset
		.in_ready          (in_ready),          //  output,    width = 1,     sink0.ready
		.in_valid          (in_valid),          //   input,    width = 1,          .valid
		.in_startofpacket  (in_startofpacket),  //   input,    width = 1,          .startofpacket
		.in_endofpacket    (in_endofpacket),    //   input,    width = 1,          .endofpacket
		.in_empty          (in_empty),          //   input,    width = 6,          .empty
		.in_error          (in_error),          //   input,    width = 1,          .error
		.in_data           (in_data),           //   input,  width = 512,          .data
		.out_ready         (out_ready),         //   input,    width = 1,   source0.ready
		.out_valid         (out_valid),         //  output,    width = 1,          .valid
		.out_startofpacket (out_startofpacket), //  output,    width = 1,          .startofpacket
		.out_endofpacket   (out_endofpacket),   //  output,    width = 1,          .endofpacket
		.out_empty         (out_empty),         //  output,    width = 6,          .empty
		.out_error         (out_error),         //  output,    width = 1,          .error
		.out_data          (out_data),          //  output,  width = 512,          .data
		.out_channel       (),                  // (terminated),                         
		.in_channel        (1'b0)               // (terminated),                         
	);

endmodule
