// Copyright (C) 2023 Intel Corporation
// SPDX-License-Identifier: MIT

`define payload_generate(PF,VF,VA) \
          local_vf_active = ``VA``;\
          local_pf_num    = ``PF``;\
          local_vf_num    = ``VF``;\
          local_tlp_length = $urandom_range(1,64) ;\
          local_payload = 'h0;\
          local_my_payload = 'h0;\
          assert(std::randomize(random_value));\      
          for(int j=0; j < (local_tlp_length*32); j++) local_my_payload[j] = 1'b1;\
          local_payload = (random_value) & local_my_payload;\
          `uvm_info("body", $sformatf("TLP Length = %h and Payload = %h and Random Value generated = %h No of Trans = %d",local_tlp_length,local_payload,random_value,no_of_transactions),UVM_LOW)\

class pf_vf_mux_stress_seq extends uvm_sequence;
    
     bit local_vf_active       ;
     bit [2:0] local_pf_num    ;
     bit [10:0] local_vf_num   ;
     bit [9:0] local_tlp_length;
     bit [255:0] local_payload , random_value, local_my_payload;
     rand int no_of_transactions ;    
     
     `ifdef TB_CONFIG_1
     int port_count[16];
     `endif
     `ifdef TB_CONFIG_2
     int port_count[24];
     `endif
     `ifdef TB_CONFIG_3
     int port_count[32];
     `endif
     `ifdef TB_CONFIG_4
     int port_count[2048];
     `endif
    
  `uvm_object_utils(pf_vf_mux_stress_seq);

  /** Declare a typed sequencer object that the sequence can access */
  `uvm_declare_p_sequencer(pf_vf_mux_virtual_sequencer)


    function new (string name = "pf_vf_mux_stress_seq");
        super.new(name);
    endfunction : new

     virtual function void build_phase(uvm_phase phase);
      endfunction: build_phase


    task body();
        pf_vf_mux_request_sequence master_seq_1,master_seq_2;
        super.body(); 
      	`uvm_info(get_name(), "Entering PF0 Traffic sequence...", UVM_LOW)
        `uvm_info(get_name(), "Starting master sequence on Host master sequencer", UVM_LOW)
        for(int i = 0; i < no_of_transactions; i++) begin
        fork
          begin 
 
              //===============================================
              // Generating the payload w.r.t TLP length field
              //===============================================
              `ifdef TB_CONFIG_1
                 local_pf_num = $urandom_range(0,7);
                 local_vf_num = 0;
                 local_vf_active = $urandom_range(0,1);
              `elsif TB_CONFIG_2
                 local_pf_num = $urandom_range(0,7);
                 if(i<(no_of_transactions/3)) begin
                   local_vf_num = 'h7FF;
                   local_vf_active = 1;
                 end
                 else begin
                   local_vf_num = 0;
                   local_vf_active = $urandom_range(0,1);
                 end
              `elsif TB_CONFIG_3
                 local_pf_num = $urandom_range(0,7);
                 if(i<=(no_of_transactions/2)) begin
                   local_vf_num = 0;
                   local_vf_active = $urandom_range(0,1);
                 end
                 else if (i<(3*(no_of_transactions/4)))begin
                   local_vf_num = 'h7FF;
                   local_vf_active = 1;
                 end
                 else begin
                   local_vf_num = `RANDOM_VF;
                   local_vf_active = 1;
                 end
               `else
                 local_pf_num = 0;
                 local_vf_num = $urandom_range(0,2047);
                 local_vf_active = 1;
               `endif
                
              local_tlp_length = $urandom_range(1,64) ;
              local_payload = 'h0;
              local_my_payload = 'h0;
              assert(std::randomize(random_value));      
             
              // For stress_test port packet count
              `ifndef TB_CONFIG_4
              if (local_pf_num == 0 && local_vf_num == 0 && local_vf_active == 0) port_count[0]++;  
              else if (local_pf_num == 1 && local_vf_num == 0 && local_vf_active == 0) port_count[1]++;  
              else if (local_pf_num == 2 && local_vf_num == 0 && local_vf_active == 0) port_count[2]++;  
              else if (local_pf_num == 3 && local_vf_num == 0 && local_vf_active == 0) port_count[3]++;  
              else if (local_pf_num == 4 && local_vf_num == 0 && local_vf_active == 0) port_count[4]++;  
              else if (local_pf_num == 5 && local_vf_num == 0 && local_vf_active == 0) port_count[5]++;  
              else if (local_pf_num == 6 && local_vf_num == 0 && local_vf_active == 0) port_count[6]++;  
              else if (local_pf_num == 7 && local_vf_num == 0 && local_vf_active == 0) port_count[7]++;  
              else if (local_pf_num == 0 && local_vf_num == 0 && local_vf_active == 1) port_count[8]++;  
              else if (local_pf_num == 1 && local_vf_num == 0 && local_vf_active == 1) port_count[9]++;  
              else if (local_pf_num == 2 && local_vf_num == 0 && local_vf_active == 1) port_count[10]++;  
              else if (local_pf_num == 3 && local_vf_num == 0 && local_vf_active == 1) port_count[11]++;  
              else if (local_pf_num == 4 && local_vf_num == 0 && local_vf_active == 1) port_count[12]++;  
              else if (local_pf_num == 5 && local_vf_num == 0 && local_vf_active == 1) port_count[13]++;  
              else if (local_pf_num == 6 && local_vf_num == 0 && local_vf_active == 1) port_count[14]++;  
              else if (local_pf_num == 7 && local_vf_num == 0 && local_vf_active == 1) port_count[15]++; 
              `ifndef TB_CONFIG_1
              else if (local_pf_num == 0 && local_vf_num == 2047 && local_vf_active == 1) port_count[16]++;  
              else if (local_pf_num == 1 && local_vf_num == 2047 && local_vf_active == 1) port_count[17]++;  
              else if (local_pf_num == 2 && local_vf_num == 2047 && local_vf_active == 1) port_count[18]++;  
              else if (local_pf_num == 3 && local_vf_num == 2047 && local_vf_active == 1) port_count[19]++;  
              else if (local_pf_num == 4 && local_vf_num == 2047 && local_vf_active == 1) port_count[20]++;  
              else if (local_pf_num == 5 && local_vf_num == 2047 && local_vf_active == 1) port_count[21]++;  
              else if (local_pf_num == 6 && local_vf_num == 2047 && local_vf_active == 1) port_count[22]++;  
              else if (local_pf_num == 7 && local_vf_num == 2047 && local_vf_active == 1) port_count[23]++;
              `endif
              `ifdef TB_CONFIG_3
              else if (local_pf_num == 0 && local_vf_num == `RANDOM_VF && local_vf_active == 1) port_count[24]++;  
              else if (local_pf_num == 1 && local_vf_num == `RANDOM_VF && local_vf_active == 1) port_count[25]++;  
              else if (local_pf_num == 2 && local_vf_num == `RANDOM_VF && local_vf_active == 1) port_count[26]++;  
              else if (local_pf_num == 3 && local_vf_num == `RANDOM_VF && local_vf_active == 1) port_count[27]++;  
              else if (local_pf_num == 4 && local_vf_num == `RANDOM_VF && local_vf_active == 1) port_count[28]++;  
              else if (local_pf_num == 5 && local_vf_num == `RANDOM_VF && local_vf_active == 1) port_count[29]++;  
              else if (local_pf_num == 6 && local_vf_num == `RANDOM_VF && local_vf_active == 1) port_count[30]++;  
              else if (local_pf_num == 7 && local_vf_num == `RANDOM_VF && local_vf_active == 1) port_count[31]++;
              `endif
              `endif
              `ifdef TB_CONFIG_4
              if (local_pf_num == 0 && local_vf_num == 0 && local_vf_active == 1) port_count[0]++;  
              else if (local_pf_num == 0 && local_vf_num == 1 && local_vf_active == 1) port_count[1]++; 
              else if (local_pf_num == 0 && local_vf_num == 2 && local_vf_active == 1) port_count[2]++; 
              else if (local_pf_num == 0 && local_vf_num == 3 && local_vf_active == 1) port_count[3]++; 
              else if (local_pf_num == 0 && local_vf_num == 4 && local_vf_active == 1) port_count[4]++; 
              else if (local_pf_num == 0 && local_vf_num == 5 && local_vf_active == 1) port_count[5]++; 
              else if (local_pf_num == 0 && local_vf_num == 6 && local_vf_active == 1) port_count[6]++; 
              else if (local_pf_num == 0 && local_vf_num == 7 && local_vf_active == 1) port_count[7]++; 
              else if (local_pf_num == 0 && local_vf_num == 8 && local_vf_active == 1) port_count[8]++; 
              else if (local_pf_num == 0 && local_vf_num == 9 && local_vf_active == 1) port_count[9]++; 
              else if (local_pf_num == 0 && local_vf_num == 10 && local_vf_active == 1) port_count[10]++; 
              else if (local_pf_num == 0 && local_vf_num == 11 && local_vf_active == 1) port_count[11]++; 
              else if (local_pf_num == 0 && local_vf_num == 12 && local_vf_active == 1) port_count[12]++; 
              else if (local_pf_num == 0 && local_vf_num == 13 && local_vf_active == 1) port_count[13]++; 
              else if (local_pf_num == 0 && local_vf_num == 14 && local_vf_active == 1) port_count[14]++; 
              else if (local_pf_num == 0 && local_vf_num == 15 && local_vf_active == 1) port_count[15]++; 
              else if (local_pf_num == 0 && local_vf_num == 16 && local_vf_active == 1) port_count[16]++; 
              else if (local_pf_num == 0 && local_vf_num == 17 && local_vf_active == 1) port_count[17]++; 
              else if (local_pf_num == 0 && local_vf_num == 18 && local_vf_active == 1) port_count[18]++; 
              else if (local_pf_num == 0 && local_vf_num == 19 && local_vf_active == 1) port_count[19]++; 
              else if (local_pf_num == 0 && local_vf_num == 20 && local_vf_active == 1) port_count[20]++; 
              else if (local_pf_num == 0 && local_vf_num == 21 && local_vf_active == 1) port_count[21]++; 
              else if (local_pf_num == 0 && local_vf_num == 22 && local_vf_active == 1) port_count[22]++; 
              else if (local_pf_num == 0 && local_vf_num == 23 && local_vf_active == 1) port_count[23]++; 
              else if (local_pf_num == 0 && local_vf_num == 24 && local_vf_active == 1) port_count[24]++; 
              else if (local_pf_num == 0 && local_vf_num == 25 && local_vf_active == 1) port_count[25]++; 
              else if (local_pf_num == 0 && local_vf_num == 26 && local_vf_active == 1) port_count[26]++; 
              else if (local_pf_num == 0 && local_vf_num == 27 && local_vf_active == 1) port_count[27]++; 
              else if (local_pf_num == 0 && local_vf_num == 28 && local_vf_active == 1) port_count[28]++; 
              else if (local_pf_num == 0 && local_vf_num == 29 && local_vf_active == 1) port_count[29]++; 
              else if (local_pf_num == 0 && local_vf_num == 30 && local_vf_active == 1) port_count[30]++; 
              else if (local_pf_num == 0 && local_vf_num == 31 && local_vf_active == 1) port_count[31]++; 
              else if (local_pf_num == 0 && local_vf_num == 32 && local_vf_active == 1) port_count[32]++; 
              else if (local_pf_num == 0 && local_vf_num == 33 && local_vf_active == 1) port_count[33]++; 
              else if (local_pf_num == 0 && local_vf_num == 34 && local_vf_active == 1) port_count[34]++; 
              else if (local_pf_num == 0 && local_vf_num == 35 && local_vf_active == 1) port_count[35]++; 
              else if (local_pf_num == 0 && local_vf_num == 36 && local_vf_active == 1) port_count[36]++; 
              else if (local_pf_num == 0 && local_vf_num == 37 && local_vf_active == 1) port_count[37]++; 
              else if (local_pf_num == 0 && local_vf_num == 38 && local_vf_active == 1) port_count[38]++; 
              else if (local_pf_num == 0 && local_vf_num == 39 && local_vf_active == 1) port_count[39]++; 
              else if (local_pf_num == 0 && local_vf_num == 40 && local_vf_active == 1) port_count[40]++; 
              else if (local_pf_num == 0 && local_vf_num == 41 && local_vf_active == 1) port_count[41]++; 
              else if (local_pf_num == 0 && local_vf_num == 42 && local_vf_active == 1) port_count[42]++; 
              else if (local_pf_num == 0 && local_vf_num == 43 && local_vf_active == 1) port_count[43]++; 
              else if (local_pf_num == 0 && local_vf_num == 44 && local_vf_active == 1) port_count[44]++; 
              else if (local_pf_num == 0 && local_vf_num == 45 && local_vf_active == 1) port_count[45]++; 
              else if (local_pf_num == 0 && local_vf_num == 46 && local_vf_active == 1) port_count[46]++; 
              else if (local_pf_num == 0 && local_vf_num == 47 && local_vf_active == 1) port_count[47]++; 
              else if (local_pf_num == 0 && local_vf_num == 48 && local_vf_active == 1) port_count[48]++; 
              else if (local_pf_num == 0 && local_vf_num == 49 && local_vf_active == 1) port_count[49]++; 
              else if (local_pf_num == 0 && local_vf_num == 50 && local_vf_active == 1) port_count[50]++; 
              else if (local_pf_num == 0 && local_vf_num == 51 && local_vf_active == 1) port_count[51]++; 
              else if (local_pf_num == 0 && local_vf_num == 52 && local_vf_active == 1) port_count[52]++; 
              else if (local_pf_num == 0 && local_vf_num == 53 && local_vf_active == 1) port_count[53]++; 
              else if (local_pf_num == 0 && local_vf_num == 54 && local_vf_active == 1) port_count[54]++; 
              else if (local_pf_num == 0 && local_vf_num == 55 && local_vf_active == 1) port_count[55]++; 
              else if (local_pf_num == 0 && local_vf_num == 56 && local_vf_active == 1) port_count[56]++; 
              else if (local_pf_num == 0 && local_vf_num == 57 && local_vf_active == 1) port_count[57]++; 
              else if (local_pf_num == 0 && local_vf_num == 58 && local_vf_active == 1) port_count[58]++; 
              else if (local_pf_num == 0 && local_vf_num == 59 && local_vf_active == 1) port_count[59]++; 
              else if (local_pf_num == 0 && local_vf_num == 60 && local_vf_active == 1) port_count[60]++; 
              else if (local_pf_num == 0 && local_vf_num == 61 && local_vf_active == 1) port_count[61]++; 
              else if (local_pf_num == 0 && local_vf_num == 62 && local_vf_active == 1) port_count[62]++; 
              else if (local_pf_num == 0 && local_vf_num == 63 && local_vf_active == 1) port_count[63]++; 
              else if (local_pf_num == 0 && local_vf_num == 64 && local_vf_active == 1) port_count[64]++; 
              else if (local_pf_num == 0 && local_vf_num == 65 && local_vf_active == 1) port_count[65]++; 
              else if (local_pf_num == 0 && local_vf_num == 66 && local_vf_active == 1) port_count[66]++; 
              else if (local_pf_num == 0 && local_vf_num == 67 && local_vf_active == 1) port_count[67]++; 
              else if (local_pf_num == 0 && local_vf_num == 68 && local_vf_active == 1) port_count[68]++; 
              else if (local_pf_num == 0 && local_vf_num == 69 && local_vf_active == 1) port_count[69]++; 
              else if (local_pf_num == 0 && local_vf_num == 70 && local_vf_active == 1) port_count[70]++; 
              else if (local_pf_num == 0 && local_vf_num == 71 && local_vf_active == 1) port_count[71]++; 
              else if (local_pf_num == 0 && local_vf_num == 72 && local_vf_active == 1) port_count[72]++; 
              else if (local_pf_num == 0 && local_vf_num == 73 && local_vf_active == 1) port_count[73]++; 
              else if (local_pf_num == 0 && local_vf_num == 74 && local_vf_active == 1) port_count[74]++; 
              else if (local_pf_num == 0 && local_vf_num == 75 && local_vf_active == 1) port_count[75]++; 
              else if (local_pf_num == 0 && local_vf_num == 76 && local_vf_active == 1) port_count[76]++; 
              else if (local_pf_num == 0 && local_vf_num == 77 && local_vf_active == 1) port_count[77]++; 
              else if (local_pf_num == 0 && local_vf_num == 78 && local_vf_active == 1) port_count[78]++; 
              else if (local_pf_num == 0 && local_vf_num == 79 && local_vf_active == 1) port_count[79]++; 
              else if (local_pf_num == 0 && local_vf_num == 80 && local_vf_active == 1) port_count[80]++; 
              else if (local_pf_num == 0 && local_vf_num == 81 && local_vf_active == 1) port_count[81]++; 
              else if (local_pf_num == 0 && local_vf_num == 82 && local_vf_active == 1) port_count[82]++; 
              else if (local_pf_num == 0 && local_vf_num == 83 && local_vf_active == 1) port_count[83]++; 
              else if (local_pf_num == 0 && local_vf_num == 84 && local_vf_active == 1) port_count[84]++; 
              else if (local_pf_num == 0 && local_vf_num == 85 && local_vf_active == 1) port_count[85]++; 
              else if (local_pf_num == 0 && local_vf_num == 86 && local_vf_active == 1) port_count[86]++; 
              else if (local_pf_num == 0 && local_vf_num == 87 && local_vf_active == 1) port_count[87]++; 
              else if (local_pf_num == 0 && local_vf_num == 88 && local_vf_active == 1) port_count[88]++; 
              else if (local_pf_num == 0 && local_vf_num == 89 && local_vf_active == 1) port_count[89]++; 
              else if (local_pf_num == 0 && local_vf_num == 90 && local_vf_active == 1) port_count[90]++; 
              else if (local_pf_num == 0 && local_vf_num == 91 && local_vf_active == 1) port_count[91]++; 
              else if (local_pf_num == 0 && local_vf_num == 92 && local_vf_active == 1) port_count[92]++; 
              else if (local_pf_num == 0 && local_vf_num == 93 && local_vf_active == 1) port_count[93]++; 
              else if (local_pf_num == 0 && local_vf_num == 94 && local_vf_active == 1) port_count[94]++; 
              else if (local_pf_num == 0 && local_vf_num == 95 && local_vf_active == 1) port_count[95]++; 
              else if (local_pf_num == 0 && local_vf_num == 96 && local_vf_active == 1) port_count[96]++; 
              else if (local_pf_num == 0 && local_vf_num == 97 && local_vf_active == 1) port_count[97]++; 
              else if (local_pf_num == 0 && local_vf_num == 98 && local_vf_active == 1) port_count[98]++; 
              else if (local_pf_num == 0 && local_vf_num == 99 && local_vf_active == 1) port_count[99]++; 
              else if (local_pf_num == 0 && local_vf_num == 100 && local_vf_active == 1) port_count[100]++; 
              else if (local_pf_num == 0 && local_vf_num == 101 && local_vf_active == 1) port_count[101]++; 
              else if (local_pf_num == 0 && local_vf_num == 102 && local_vf_active == 1) port_count[102]++; 
              else if (local_pf_num == 0 && local_vf_num == 103 && local_vf_active == 1) port_count[103]++; 
              else if (local_pf_num == 0 && local_vf_num == 104 && local_vf_active == 1) port_count[104]++; 
              else if (local_pf_num == 0 && local_vf_num == 105 && local_vf_active == 1) port_count[105]++; 
              else if (local_pf_num == 0 && local_vf_num == 106 && local_vf_active == 1) port_count[106]++; 
              else if (local_pf_num == 0 && local_vf_num == 107 && local_vf_active == 1) port_count[107]++; 
              else if (local_pf_num == 0 && local_vf_num == 108 && local_vf_active == 1) port_count[108]++; 
              else if (local_pf_num == 0 && local_vf_num == 109 && local_vf_active == 1) port_count[109]++; 
              else if (local_pf_num == 0 && local_vf_num == 110 && local_vf_active == 1) port_count[110]++; 
              else if (local_pf_num == 0 && local_vf_num == 111 && local_vf_active == 1) port_count[111]++; 
              else if (local_pf_num == 0 && local_vf_num == 112 && local_vf_active == 1) port_count[112]++; 
              else if (local_pf_num == 0 && local_vf_num == 113 && local_vf_active == 1) port_count[113]++; 
              else if (local_pf_num == 0 && local_vf_num == 114 && local_vf_active == 1) port_count[114]++; 
              else if (local_pf_num == 0 && local_vf_num == 115 && local_vf_active == 1) port_count[115]++; 
              else if (local_pf_num == 0 && local_vf_num == 116 && local_vf_active == 1) port_count[116]++; 
              else if (local_pf_num == 0 && local_vf_num == 117 && local_vf_active == 1) port_count[117]++; 
              else if (local_pf_num == 0 && local_vf_num == 118 && local_vf_active == 1) port_count[118]++; 
              else if (local_pf_num == 0 && local_vf_num == 119 && local_vf_active == 1) port_count[119]++; 
              else if (local_pf_num == 0 && local_vf_num == 120 && local_vf_active == 1) port_count[120]++; 
              else if (local_pf_num == 0 && local_vf_num == 121 && local_vf_active == 1) port_count[121]++; 
              else if (local_pf_num == 0 && local_vf_num == 122 && local_vf_active == 1) port_count[122]++; 
              else if (local_pf_num == 0 && local_vf_num == 123 && local_vf_active == 1) port_count[123]++; 
              else if (local_pf_num == 0 && local_vf_num == 124 && local_vf_active == 1) port_count[124]++; 
              else if (local_pf_num == 0 && local_vf_num == 125 && local_vf_active == 1) port_count[125]++; 
              else if (local_pf_num == 0 && local_vf_num == 126 && local_vf_active == 1) port_count[126]++; 
              else if (local_pf_num == 0 && local_vf_num == 127 && local_vf_active == 1) port_count[127]++; 
              else if (local_pf_num == 0 && local_vf_num == 128 && local_vf_active == 1) port_count[128]++; 
              else if (local_pf_num == 0 && local_vf_num == 129 && local_vf_active == 1) port_count[129]++; 
              else if (local_pf_num == 0 && local_vf_num == 130 && local_vf_active == 1) port_count[130]++; 
              else if (local_pf_num == 0 && local_vf_num == 131 && local_vf_active == 1) port_count[131]++; 
              else if (local_pf_num == 0 && local_vf_num == 132 && local_vf_active == 1) port_count[132]++; 
              else if (local_pf_num == 0 && local_vf_num == 133 && local_vf_active == 1) port_count[133]++; 
              else if (local_pf_num == 0 && local_vf_num == 134 && local_vf_active == 1) port_count[134]++; 
              else if (local_pf_num == 0 && local_vf_num == 135 && local_vf_active == 1) port_count[135]++; 
              else if (local_pf_num == 0 && local_vf_num == 136 && local_vf_active == 1) port_count[136]++; 
              else if (local_pf_num == 0 && local_vf_num == 137 && local_vf_active == 1) port_count[137]++; 
              else if (local_pf_num == 0 && local_vf_num == 138 && local_vf_active == 1) port_count[138]++; 
              else if (local_pf_num == 0 && local_vf_num == 139 && local_vf_active == 1) port_count[139]++; 
              else if (local_pf_num == 0 && local_vf_num == 140 && local_vf_active == 1) port_count[140]++; 
              else if (local_pf_num == 0 && local_vf_num == 141 && local_vf_active == 1) port_count[141]++; 
              else if (local_pf_num == 0 && local_vf_num == 142 && local_vf_active == 1) port_count[142]++; 
              else if (local_pf_num == 0 && local_vf_num == 143 && local_vf_active == 1) port_count[143]++; 
              else if (local_pf_num == 0 && local_vf_num == 144 && local_vf_active == 1) port_count[144]++; 
              else if (local_pf_num == 0 && local_vf_num == 145 && local_vf_active == 1) port_count[145]++; 
              else if (local_pf_num == 0 && local_vf_num == 146 && local_vf_active == 1) port_count[146]++; 
              else if (local_pf_num == 0 && local_vf_num == 147 && local_vf_active == 1) port_count[147]++; 
              else if (local_pf_num == 0 && local_vf_num == 148 && local_vf_active == 1) port_count[148]++; 
              else if (local_pf_num == 0 && local_vf_num == 149 && local_vf_active == 1) port_count[149]++; 
              else if (local_pf_num == 0 && local_vf_num == 150 && local_vf_active == 1) port_count[150]++; 
              else if (local_pf_num == 0 && local_vf_num == 151 && local_vf_active == 1) port_count[151]++; 
              else if (local_pf_num == 0 && local_vf_num == 152 && local_vf_active == 1) port_count[152]++; 
              else if (local_pf_num == 0 && local_vf_num == 153 && local_vf_active == 1) port_count[153]++; 
              else if (local_pf_num == 0 && local_vf_num == 154 && local_vf_active == 1) port_count[154]++; 
              else if (local_pf_num == 0 && local_vf_num == 155 && local_vf_active == 1) port_count[155]++; 
              else if (local_pf_num == 0 && local_vf_num == 156 && local_vf_active == 1) port_count[156]++; 
              else if (local_pf_num == 0 && local_vf_num == 157 && local_vf_active == 1) port_count[157]++; 
              else if (local_pf_num == 0 && local_vf_num == 158 && local_vf_active == 1) port_count[158]++; 
              else if (local_pf_num == 0 && local_vf_num == 159 && local_vf_active == 1) port_count[159]++; 
              else if (local_pf_num == 0 && local_vf_num == 160 && local_vf_active == 1) port_count[160]++; 
              else if (local_pf_num == 0 && local_vf_num == 161 && local_vf_active == 1) port_count[161]++; 
              else if (local_pf_num == 0 && local_vf_num == 162 && local_vf_active == 1) port_count[162]++; 
              else if (local_pf_num == 0 && local_vf_num == 163 && local_vf_active == 1) port_count[163]++; 
              else if (local_pf_num == 0 && local_vf_num == 164 && local_vf_active == 1) port_count[164]++; 
              else if (local_pf_num == 0 && local_vf_num == 165 && local_vf_active == 1) port_count[165]++; 
              else if (local_pf_num == 0 && local_vf_num == 166 && local_vf_active == 1) port_count[166]++; 
              else if (local_pf_num == 0 && local_vf_num == 167 && local_vf_active == 1) port_count[167]++; 
              else if (local_pf_num == 0 && local_vf_num == 168 && local_vf_active == 1) port_count[168]++; 
              else if (local_pf_num == 0 && local_vf_num == 169 && local_vf_active == 1) port_count[169]++; 
              else if (local_pf_num == 0 && local_vf_num == 170 && local_vf_active == 1) port_count[170]++; 
              else if (local_pf_num == 0 && local_vf_num == 171 && local_vf_active == 1) port_count[171]++; 
              else if (local_pf_num == 0 && local_vf_num == 172 && local_vf_active == 1) port_count[172]++; 
              else if (local_pf_num == 0 && local_vf_num == 173 && local_vf_active == 1) port_count[173]++; 
              else if (local_pf_num == 0 && local_vf_num == 174 && local_vf_active == 1) port_count[174]++; 
              else if (local_pf_num == 0 && local_vf_num == 175 && local_vf_active == 1) port_count[175]++; 
              else if (local_pf_num == 0 && local_vf_num == 176 && local_vf_active == 1) port_count[176]++; 
              else if (local_pf_num == 0 && local_vf_num == 177 && local_vf_active == 1) port_count[177]++; 
              else if (local_pf_num == 0 && local_vf_num == 178 && local_vf_active == 1) port_count[178]++; 
              else if (local_pf_num == 0 && local_vf_num == 179 && local_vf_active == 1) port_count[179]++; 
              else if (local_pf_num == 0 && local_vf_num == 180 && local_vf_active == 1) port_count[180]++; 
              else if (local_pf_num == 0 && local_vf_num == 181 && local_vf_active == 1) port_count[181]++; 
              else if (local_pf_num == 0 && local_vf_num == 182 && local_vf_active == 1) port_count[182]++; 
              else if (local_pf_num == 0 && local_vf_num == 183 && local_vf_active == 1) port_count[183]++; 
              else if (local_pf_num == 0 && local_vf_num == 184 && local_vf_active == 1) port_count[184]++; 
              else if (local_pf_num == 0 && local_vf_num == 185 && local_vf_active == 1) port_count[185]++; 
              else if (local_pf_num == 0 && local_vf_num == 186 && local_vf_active == 1) port_count[186]++; 
              else if (local_pf_num == 0 && local_vf_num == 187 && local_vf_active == 1) port_count[187]++; 
              else if (local_pf_num == 0 && local_vf_num == 188 && local_vf_active == 1) port_count[188]++; 
              else if (local_pf_num == 0 && local_vf_num == 189 && local_vf_active == 1) port_count[189]++; 
              else if (local_pf_num == 0 && local_vf_num == 190 && local_vf_active == 1) port_count[190]++; 
              else if (local_pf_num == 0 && local_vf_num == 191 && local_vf_active == 1) port_count[191]++; 
              else if (local_pf_num == 0 && local_vf_num == 192 && local_vf_active == 1) port_count[192]++; 
              else if (local_pf_num == 0 && local_vf_num == 193 && local_vf_active == 1) port_count[193]++; 
              else if (local_pf_num == 0 && local_vf_num == 194 && local_vf_active == 1) port_count[194]++; 
              else if (local_pf_num == 0 && local_vf_num == 195 && local_vf_active == 1) port_count[195]++; 
              else if (local_pf_num == 0 && local_vf_num == 196 && local_vf_active == 1) port_count[196]++; 
              else if (local_pf_num == 0 && local_vf_num == 197 && local_vf_active == 1) port_count[197]++; 
              else if (local_pf_num == 0 && local_vf_num == 198 && local_vf_active == 1) port_count[198]++; 
              else if (local_pf_num == 0 && local_vf_num == 199 && local_vf_active == 1) port_count[199]++; 
              else if (local_pf_num == 0 && local_vf_num == 200 && local_vf_active == 1) port_count[200]++; 
              else if (local_pf_num == 0 && local_vf_num == 201 && local_vf_active == 1) port_count[201]++; 
              else if (local_pf_num == 0 && local_vf_num == 202 && local_vf_active == 1) port_count[202]++; 
              else if (local_pf_num == 0 && local_vf_num == 203 && local_vf_active == 1) port_count[203]++; 
              else if (local_pf_num == 0 && local_vf_num == 204 && local_vf_active == 1) port_count[204]++; 
              else if (local_pf_num == 0 && local_vf_num == 205 && local_vf_active == 1) port_count[205]++; 
              else if (local_pf_num == 0 && local_vf_num == 206 && local_vf_active == 1) port_count[206]++; 
              else if (local_pf_num == 0 && local_vf_num == 207 && local_vf_active == 1) port_count[207]++; 
              else if (local_pf_num == 0 && local_vf_num == 208 && local_vf_active == 1) port_count[208]++; 
              else if (local_pf_num == 0 && local_vf_num == 209 && local_vf_active == 1) port_count[209]++; 
              else if (local_pf_num == 0 && local_vf_num == 210 && local_vf_active == 1) port_count[210]++; 
              else if (local_pf_num == 0 && local_vf_num == 211 && local_vf_active == 1) port_count[211]++; 
              else if (local_pf_num == 0 && local_vf_num == 212 && local_vf_active == 1) port_count[212]++; 
              else if (local_pf_num == 0 && local_vf_num == 213 && local_vf_active == 1) port_count[213]++; 
              else if (local_pf_num == 0 && local_vf_num == 214 && local_vf_active == 1) port_count[214]++; 
              else if (local_pf_num == 0 && local_vf_num == 215 && local_vf_active == 1) port_count[215]++; 
              else if (local_pf_num == 0 && local_vf_num == 216 && local_vf_active == 1) port_count[216]++; 
              else if (local_pf_num == 0 && local_vf_num == 217 && local_vf_active == 1) port_count[217]++; 
              else if (local_pf_num == 0 && local_vf_num == 218 && local_vf_active == 1) port_count[218]++; 
              else if (local_pf_num == 0 && local_vf_num == 219 && local_vf_active == 1) port_count[219]++; 
              else if (local_pf_num == 0 && local_vf_num == 220 && local_vf_active == 1) port_count[220]++; 
              else if (local_pf_num == 0 && local_vf_num == 221 && local_vf_active == 1) port_count[221]++; 
              else if (local_pf_num == 0 && local_vf_num == 222 && local_vf_active == 1) port_count[222]++; 
              else if (local_pf_num == 0 && local_vf_num == 223 && local_vf_active == 1) port_count[223]++; 
              else if (local_pf_num == 0 && local_vf_num == 224 && local_vf_active == 1) port_count[224]++; 
              else if (local_pf_num == 0 && local_vf_num == 225 && local_vf_active == 1) port_count[225]++; 
              else if (local_pf_num == 0 && local_vf_num == 226 && local_vf_active == 1) port_count[226]++; 
              else if (local_pf_num == 0 && local_vf_num == 227 && local_vf_active == 1) port_count[227]++; 
              else if (local_pf_num == 0 && local_vf_num == 228 && local_vf_active == 1) port_count[228]++; 
              else if (local_pf_num == 0 && local_vf_num == 229 && local_vf_active == 1) port_count[229]++; 
              else if (local_pf_num == 0 && local_vf_num == 230 && local_vf_active == 1) port_count[230]++; 
              else if (local_pf_num == 0 && local_vf_num == 231 && local_vf_active == 1) port_count[231]++; 
              else if (local_pf_num == 0 && local_vf_num == 232 && local_vf_active == 1) port_count[232]++; 
              else if (local_pf_num == 0 && local_vf_num == 233 && local_vf_active == 1) port_count[233]++; 
              else if (local_pf_num == 0 && local_vf_num == 234 && local_vf_active == 1) port_count[234]++; 
              else if (local_pf_num == 0 && local_vf_num == 235 && local_vf_active == 1) port_count[235]++; 
              else if (local_pf_num == 0 && local_vf_num == 236 && local_vf_active == 1) port_count[236]++; 
              else if (local_pf_num == 0 && local_vf_num == 237 && local_vf_active == 1) port_count[237]++; 
              else if (local_pf_num == 0 && local_vf_num == 238 && local_vf_active == 1) port_count[238]++; 
              else if (local_pf_num == 0 && local_vf_num == 239 && local_vf_active == 1) port_count[239]++; 
              else if (local_pf_num == 0 && local_vf_num == 240 && local_vf_active == 1) port_count[240]++; 
              else if (local_pf_num == 0 && local_vf_num == 241 && local_vf_active == 1) port_count[241]++; 
              else if (local_pf_num == 0 && local_vf_num == 242 && local_vf_active == 1) port_count[242]++; 
              else if (local_pf_num == 0 && local_vf_num == 243 && local_vf_active == 1) port_count[243]++; 
              else if (local_pf_num == 0 && local_vf_num == 244 && local_vf_active == 1) port_count[244]++; 
              else if (local_pf_num == 0 && local_vf_num == 245 && local_vf_active == 1) port_count[245]++; 
              else if (local_pf_num == 0 && local_vf_num == 246 && local_vf_active == 1) port_count[246]++; 
              else if (local_pf_num == 0 && local_vf_num == 247 && local_vf_active == 1) port_count[247]++; 
              else if (local_pf_num == 0 && local_vf_num == 248 && local_vf_active == 1) port_count[248]++; 
              else if (local_pf_num == 0 && local_vf_num == 249 && local_vf_active == 1) port_count[249]++; 
              else if (local_pf_num == 0 && local_vf_num == 250 && local_vf_active == 1) port_count[250]++; 
              else if (local_pf_num == 0 && local_vf_num == 251 && local_vf_active == 1) port_count[251]++; 
              else if (local_pf_num == 0 && local_vf_num == 252 && local_vf_active == 1) port_count[252]++; 
              else if (local_pf_num == 0 && local_vf_num == 253 && local_vf_active == 1) port_count[253]++; 
              else if (local_pf_num == 0 && local_vf_num == 254 && local_vf_active == 1) port_count[254]++; 
              else if (local_pf_num == 0 && local_vf_num == 255 && local_vf_active == 1) port_count[255]++; 
              else if (local_pf_num == 0 && local_vf_num == 256 && local_vf_active == 1) port_count[256]++; 
              else if (local_pf_num == 0 && local_vf_num == 257 && local_vf_active == 1) port_count[257]++; 
              else if (local_pf_num == 0 && local_vf_num == 258 && local_vf_active == 1) port_count[258]++; 
              else if (local_pf_num == 0 && local_vf_num == 259 && local_vf_active == 1) port_count[259]++; 
              else if (local_pf_num == 0 && local_vf_num == 260 && local_vf_active == 1) port_count[260]++; 
              else if (local_pf_num == 0 && local_vf_num == 261 && local_vf_active == 1) port_count[261]++; 
              else if (local_pf_num == 0 && local_vf_num == 262 && local_vf_active == 1) port_count[262]++; 
              else if (local_pf_num == 0 && local_vf_num == 263 && local_vf_active == 1) port_count[263]++; 
              else if (local_pf_num == 0 && local_vf_num == 264 && local_vf_active == 1) port_count[264]++; 
              else if (local_pf_num == 0 && local_vf_num == 265 && local_vf_active == 1) port_count[265]++; 
              else if (local_pf_num == 0 && local_vf_num == 266 && local_vf_active == 1) port_count[266]++; 
              else if (local_pf_num == 0 && local_vf_num == 267 && local_vf_active == 1) port_count[267]++; 
              else if (local_pf_num == 0 && local_vf_num == 268 && local_vf_active == 1) port_count[268]++; 
              else if (local_pf_num == 0 && local_vf_num == 269 && local_vf_active == 1) port_count[269]++; 
              else if (local_pf_num == 0 && local_vf_num == 270 && local_vf_active == 1) port_count[270]++; 
              else if (local_pf_num == 0 && local_vf_num == 271 && local_vf_active == 1) port_count[271]++; 
              else if (local_pf_num == 0 && local_vf_num == 272 && local_vf_active == 1) port_count[272]++; 
              else if (local_pf_num == 0 && local_vf_num == 273 && local_vf_active == 1) port_count[273]++; 
              else if (local_pf_num == 0 && local_vf_num == 274 && local_vf_active == 1) port_count[274]++; 
              else if (local_pf_num == 0 && local_vf_num == 275 && local_vf_active == 1) port_count[275]++; 
              else if (local_pf_num == 0 && local_vf_num == 276 && local_vf_active == 1) port_count[276]++; 
              else if (local_pf_num == 0 && local_vf_num == 277 && local_vf_active == 1) port_count[277]++; 
              else if (local_pf_num == 0 && local_vf_num == 278 && local_vf_active == 1) port_count[278]++; 
              else if (local_pf_num == 0 && local_vf_num == 279 && local_vf_active == 1) port_count[279]++; 
              else if (local_pf_num == 0 && local_vf_num == 280 && local_vf_active == 1) port_count[280]++; 
              else if (local_pf_num == 0 && local_vf_num == 281 && local_vf_active == 1) port_count[281]++; 
              else if (local_pf_num == 0 && local_vf_num == 282 && local_vf_active == 1) port_count[282]++; 
              else if (local_pf_num == 0 && local_vf_num == 283 && local_vf_active == 1) port_count[283]++; 
              else if (local_pf_num == 0 && local_vf_num == 284 && local_vf_active == 1) port_count[284]++; 
              else if (local_pf_num == 0 && local_vf_num == 285 && local_vf_active == 1) port_count[285]++; 
              else if (local_pf_num == 0 && local_vf_num == 286 && local_vf_active == 1) port_count[286]++; 
              else if (local_pf_num == 0 && local_vf_num == 287 && local_vf_active == 1) port_count[287]++; 
              else if (local_pf_num == 0 && local_vf_num == 288 && local_vf_active == 1) port_count[288]++; 
              else if (local_pf_num == 0 && local_vf_num == 289 && local_vf_active == 1) port_count[289]++; 
              else if (local_pf_num == 0 && local_vf_num == 290 && local_vf_active == 1) port_count[290]++; 
              else if (local_pf_num == 0 && local_vf_num == 291 && local_vf_active == 1) port_count[291]++; 
              else if (local_pf_num == 0 && local_vf_num == 292 && local_vf_active == 1) port_count[292]++; 
              else if (local_pf_num == 0 && local_vf_num == 293 && local_vf_active == 1) port_count[293]++; 
              else if (local_pf_num == 0 && local_vf_num == 294 && local_vf_active == 1) port_count[294]++; 
              else if (local_pf_num == 0 && local_vf_num == 295 && local_vf_active == 1) port_count[295]++; 
              else if (local_pf_num == 0 && local_vf_num == 296 && local_vf_active == 1) port_count[296]++; 
              else if (local_pf_num == 0 && local_vf_num == 297 && local_vf_active == 1) port_count[297]++; 
              else if (local_pf_num == 0 && local_vf_num == 298 && local_vf_active == 1) port_count[298]++; 
              else if (local_pf_num == 0 && local_vf_num == 299 && local_vf_active == 1) port_count[299]++; 
              else if (local_pf_num == 0 && local_vf_num == 300 && local_vf_active == 1) port_count[300]++; 
              else if (local_pf_num == 0 && local_vf_num == 301 && local_vf_active == 1) port_count[301]++; 
              else if (local_pf_num == 0 && local_vf_num == 302 && local_vf_active == 1) port_count[302]++; 
              else if (local_pf_num == 0 && local_vf_num == 303 && local_vf_active == 1) port_count[303]++; 
              else if (local_pf_num == 0 && local_vf_num == 304 && local_vf_active == 1) port_count[304]++; 
              else if (local_pf_num == 0 && local_vf_num == 305 && local_vf_active == 1) port_count[305]++; 
              else if (local_pf_num == 0 && local_vf_num == 306 && local_vf_active == 1) port_count[306]++; 
              else if (local_pf_num == 0 && local_vf_num == 307 && local_vf_active == 1) port_count[307]++; 
              else if (local_pf_num == 0 && local_vf_num == 308 && local_vf_active == 1) port_count[308]++; 
              else if (local_pf_num == 0 && local_vf_num == 309 && local_vf_active == 1) port_count[309]++; 
              else if (local_pf_num == 0 && local_vf_num == 310 && local_vf_active == 1) port_count[310]++; 
              else if (local_pf_num == 0 && local_vf_num == 311 && local_vf_active == 1) port_count[311]++; 
              else if (local_pf_num == 0 && local_vf_num == 312 && local_vf_active == 1) port_count[312]++; 
              else if (local_pf_num == 0 && local_vf_num == 313 && local_vf_active == 1) port_count[313]++; 
              else if (local_pf_num == 0 && local_vf_num == 314 && local_vf_active == 1) port_count[314]++; 
              else if (local_pf_num == 0 && local_vf_num == 315 && local_vf_active == 1) port_count[315]++; 
              else if (local_pf_num == 0 && local_vf_num == 316 && local_vf_active == 1) port_count[316]++; 
              else if (local_pf_num == 0 && local_vf_num == 317 && local_vf_active == 1) port_count[317]++; 
              else if (local_pf_num == 0 && local_vf_num == 318 && local_vf_active == 1) port_count[318]++; 
              else if (local_pf_num == 0 && local_vf_num == 319 && local_vf_active == 1) port_count[319]++; 
              else if (local_pf_num == 0 && local_vf_num == 320 && local_vf_active == 1) port_count[320]++; 
              else if (local_pf_num == 0 && local_vf_num == 321 && local_vf_active == 1) port_count[321]++; 
              else if (local_pf_num == 0 && local_vf_num == 322 && local_vf_active == 1) port_count[322]++; 
              else if (local_pf_num == 0 && local_vf_num == 323 && local_vf_active == 1) port_count[323]++; 
              else if (local_pf_num == 0 && local_vf_num == 324 && local_vf_active == 1) port_count[324]++; 
              else if (local_pf_num == 0 && local_vf_num == 325 && local_vf_active == 1) port_count[325]++; 
              else if (local_pf_num == 0 && local_vf_num == 326 && local_vf_active == 1) port_count[326]++; 
              else if (local_pf_num == 0 && local_vf_num == 327 && local_vf_active == 1) port_count[327]++; 
              else if (local_pf_num == 0 && local_vf_num == 328 && local_vf_active == 1) port_count[328]++; 
              else if (local_pf_num == 0 && local_vf_num == 329 && local_vf_active == 1) port_count[329]++; 
              else if (local_pf_num == 0 && local_vf_num == 330 && local_vf_active == 1) port_count[330]++; 
              else if (local_pf_num == 0 && local_vf_num == 331 && local_vf_active == 1) port_count[331]++; 
              else if (local_pf_num == 0 && local_vf_num == 332 && local_vf_active == 1) port_count[332]++; 
              else if (local_pf_num == 0 && local_vf_num == 333 && local_vf_active == 1) port_count[333]++; 
              else if (local_pf_num == 0 && local_vf_num == 334 && local_vf_active == 1) port_count[334]++; 
              else if (local_pf_num == 0 && local_vf_num == 335 && local_vf_active == 1) port_count[335]++; 
              else if (local_pf_num == 0 && local_vf_num == 336 && local_vf_active == 1) port_count[336]++; 
              else if (local_pf_num == 0 && local_vf_num == 337 && local_vf_active == 1) port_count[337]++; 
              else if (local_pf_num == 0 && local_vf_num == 338 && local_vf_active == 1) port_count[338]++; 
              else if (local_pf_num == 0 && local_vf_num == 339 && local_vf_active == 1) port_count[339]++; 
              else if (local_pf_num == 0 && local_vf_num == 340 && local_vf_active == 1) port_count[340]++; 
              else if (local_pf_num == 0 && local_vf_num == 341 && local_vf_active == 1) port_count[341]++; 
              else if (local_pf_num == 0 && local_vf_num == 342 && local_vf_active == 1) port_count[342]++; 
              else if (local_pf_num == 0 && local_vf_num == 343 && local_vf_active == 1) port_count[343]++; 
              else if (local_pf_num == 0 && local_vf_num == 344 && local_vf_active == 1) port_count[344]++; 
              else if (local_pf_num == 0 && local_vf_num == 345 && local_vf_active == 1) port_count[345]++; 
              else if (local_pf_num == 0 && local_vf_num == 346 && local_vf_active == 1) port_count[346]++; 
              else if (local_pf_num == 0 && local_vf_num == 347 && local_vf_active == 1) port_count[347]++; 
              else if (local_pf_num == 0 && local_vf_num == 348 && local_vf_active == 1) port_count[348]++; 
              else if (local_pf_num == 0 && local_vf_num == 349 && local_vf_active == 1) port_count[349]++; 
              else if (local_pf_num == 0 && local_vf_num == 350 && local_vf_active == 1) port_count[350]++; 
              else if (local_pf_num == 0 && local_vf_num == 351 && local_vf_active == 1) port_count[351]++; 
              else if (local_pf_num == 0 && local_vf_num == 352 && local_vf_active == 1) port_count[352]++; 
              else if (local_pf_num == 0 && local_vf_num == 353 && local_vf_active == 1) port_count[353]++; 
              else if (local_pf_num == 0 && local_vf_num == 354 && local_vf_active == 1) port_count[354]++; 
              else if (local_pf_num == 0 && local_vf_num == 355 && local_vf_active == 1) port_count[355]++; 
              else if (local_pf_num == 0 && local_vf_num == 356 && local_vf_active == 1) port_count[356]++; 
              else if (local_pf_num == 0 && local_vf_num == 357 && local_vf_active == 1) port_count[357]++; 
              else if (local_pf_num == 0 && local_vf_num == 358 && local_vf_active == 1) port_count[358]++; 
              else if (local_pf_num == 0 && local_vf_num == 359 && local_vf_active == 1) port_count[359]++; 
              else if (local_pf_num == 0 && local_vf_num == 360 && local_vf_active == 1) port_count[360]++; 
              else if (local_pf_num == 0 && local_vf_num == 361 && local_vf_active == 1) port_count[361]++; 
              else if (local_pf_num == 0 && local_vf_num == 362 && local_vf_active == 1) port_count[362]++; 
              else if (local_pf_num == 0 && local_vf_num == 363 && local_vf_active == 1) port_count[363]++; 
              else if (local_pf_num == 0 && local_vf_num == 364 && local_vf_active == 1) port_count[364]++; 
              else if (local_pf_num == 0 && local_vf_num == 365 && local_vf_active == 1) port_count[365]++; 
              else if (local_pf_num == 0 && local_vf_num == 366 && local_vf_active == 1) port_count[366]++; 
              else if (local_pf_num == 0 && local_vf_num == 367 && local_vf_active == 1) port_count[367]++; 
              else if (local_pf_num == 0 && local_vf_num == 368 && local_vf_active == 1) port_count[368]++; 
              else if (local_pf_num == 0 && local_vf_num == 369 && local_vf_active == 1) port_count[369]++; 
              else if (local_pf_num == 0 && local_vf_num == 370 && local_vf_active == 1) port_count[370]++; 
              else if (local_pf_num == 0 && local_vf_num == 371 && local_vf_active == 1) port_count[371]++; 
              else if (local_pf_num == 0 && local_vf_num == 372 && local_vf_active == 1) port_count[372]++; 
              else if (local_pf_num == 0 && local_vf_num == 373 && local_vf_active == 1) port_count[373]++; 
              else if (local_pf_num == 0 && local_vf_num == 374 && local_vf_active == 1) port_count[374]++; 
              else if (local_pf_num == 0 && local_vf_num == 375 && local_vf_active == 1) port_count[375]++; 
              else if (local_pf_num == 0 && local_vf_num == 376 && local_vf_active == 1) port_count[376]++; 
              else if (local_pf_num == 0 && local_vf_num == 377 && local_vf_active == 1) port_count[377]++; 
              else if (local_pf_num == 0 && local_vf_num == 378 && local_vf_active == 1) port_count[378]++; 
              else if (local_pf_num == 0 && local_vf_num == 379 && local_vf_active == 1) port_count[379]++; 
              else if (local_pf_num == 0 && local_vf_num == 380 && local_vf_active == 1) port_count[380]++; 
              else if (local_pf_num == 0 && local_vf_num == 381 && local_vf_active == 1) port_count[381]++; 
              else if (local_pf_num == 0 && local_vf_num == 382 && local_vf_active == 1) port_count[382]++; 
              else if (local_pf_num == 0 && local_vf_num == 383 && local_vf_active == 1) port_count[383]++; 
              else if (local_pf_num == 0 && local_vf_num == 384 && local_vf_active == 1) port_count[384]++; 
              else if (local_pf_num == 0 && local_vf_num == 385 && local_vf_active == 1) port_count[385]++; 
              else if (local_pf_num == 0 && local_vf_num == 386 && local_vf_active == 1) port_count[386]++; 
              else if (local_pf_num == 0 && local_vf_num == 387 && local_vf_active == 1) port_count[387]++; 
              else if (local_pf_num == 0 && local_vf_num == 388 && local_vf_active == 1) port_count[388]++; 
              else if (local_pf_num == 0 && local_vf_num == 389 && local_vf_active == 1) port_count[389]++; 
              else if (local_pf_num == 0 && local_vf_num == 390 && local_vf_active == 1) port_count[390]++; 
              else if (local_pf_num == 0 && local_vf_num == 391 && local_vf_active == 1) port_count[391]++; 
              else if (local_pf_num == 0 && local_vf_num == 392 && local_vf_active == 1) port_count[392]++; 
              else if (local_pf_num == 0 && local_vf_num == 393 && local_vf_active == 1) port_count[393]++; 
              else if (local_pf_num == 0 && local_vf_num == 394 && local_vf_active == 1) port_count[394]++; 
              else if (local_pf_num == 0 && local_vf_num == 395 && local_vf_active == 1) port_count[395]++; 
              else if (local_pf_num == 0 && local_vf_num == 396 && local_vf_active == 1) port_count[396]++; 
              else if (local_pf_num == 0 && local_vf_num == 397 && local_vf_active == 1) port_count[397]++; 
              else if (local_pf_num == 0 && local_vf_num == 398 && local_vf_active == 1) port_count[398]++; 
              else if (local_pf_num == 0 && local_vf_num == 399 && local_vf_active == 1) port_count[399]++; 
              else if (local_pf_num == 0 && local_vf_num == 400 && local_vf_active == 1) port_count[400]++; 
              else if (local_pf_num == 0 && local_vf_num == 401 && local_vf_active == 1) port_count[401]++; 
              else if (local_pf_num == 0 && local_vf_num == 402 && local_vf_active == 1) port_count[402]++; 
              else if (local_pf_num == 0 && local_vf_num == 403 && local_vf_active == 1) port_count[403]++; 
              else if (local_pf_num == 0 && local_vf_num == 404 && local_vf_active == 1) port_count[404]++; 
              else if (local_pf_num == 0 && local_vf_num == 405 && local_vf_active == 1) port_count[405]++; 
              else if (local_pf_num == 0 && local_vf_num == 406 && local_vf_active == 1) port_count[406]++; 
              else if (local_pf_num == 0 && local_vf_num == 407 && local_vf_active == 1) port_count[407]++; 
              else if (local_pf_num == 0 && local_vf_num == 408 && local_vf_active == 1) port_count[408]++; 
              else if (local_pf_num == 0 && local_vf_num == 409 && local_vf_active == 1) port_count[409]++; 
              else if (local_pf_num == 0 && local_vf_num == 410 && local_vf_active == 1) port_count[410]++; 
              else if (local_pf_num == 0 && local_vf_num == 411 && local_vf_active == 1) port_count[411]++; 
              else if (local_pf_num == 0 && local_vf_num == 412 && local_vf_active == 1) port_count[412]++; 
              else if (local_pf_num == 0 && local_vf_num == 413 && local_vf_active == 1) port_count[413]++; 
              else if (local_pf_num == 0 && local_vf_num == 414 && local_vf_active == 1) port_count[414]++; 
              else if (local_pf_num == 0 && local_vf_num == 415 && local_vf_active == 1) port_count[415]++; 
              else if (local_pf_num == 0 && local_vf_num == 416 && local_vf_active == 1) port_count[416]++; 
              else if (local_pf_num == 0 && local_vf_num == 417 && local_vf_active == 1) port_count[417]++; 
              else if (local_pf_num == 0 && local_vf_num == 418 && local_vf_active == 1) port_count[418]++; 
              else if (local_pf_num == 0 && local_vf_num == 419 && local_vf_active == 1) port_count[419]++; 
              else if (local_pf_num == 0 && local_vf_num == 420 && local_vf_active == 1) port_count[420]++; 
              else if (local_pf_num == 0 && local_vf_num == 421 && local_vf_active == 1) port_count[421]++; 
              else if (local_pf_num == 0 && local_vf_num == 422 && local_vf_active == 1) port_count[422]++; 
              else if (local_pf_num == 0 && local_vf_num == 423 && local_vf_active == 1) port_count[423]++; 
              else if (local_pf_num == 0 && local_vf_num == 424 && local_vf_active == 1) port_count[424]++; 
              else if (local_pf_num == 0 && local_vf_num == 425 && local_vf_active == 1) port_count[425]++; 
              else if (local_pf_num == 0 && local_vf_num == 426 && local_vf_active == 1) port_count[426]++; 
              else if (local_pf_num == 0 && local_vf_num == 427 && local_vf_active == 1) port_count[427]++; 
              else if (local_pf_num == 0 && local_vf_num == 428 && local_vf_active == 1) port_count[428]++; 
              else if (local_pf_num == 0 && local_vf_num == 429 && local_vf_active == 1) port_count[429]++; 
              else if (local_pf_num == 0 && local_vf_num == 430 && local_vf_active == 1) port_count[430]++; 
              else if (local_pf_num == 0 && local_vf_num == 431 && local_vf_active == 1) port_count[431]++; 
              else if (local_pf_num == 0 && local_vf_num == 432 && local_vf_active == 1) port_count[432]++; 
              else if (local_pf_num == 0 && local_vf_num == 433 && local_vf_active == 1) port_count[433]++; 
              else if (local_pf_num == 0 && local_vf_num == 434 && local_vf_active == 1) port_count[434]++; 
              else if (local_pf_num == 0 && local_vf_num == 435 && local_vf_active == 1) port_count[435]++; 
              else if (local_pf_num == 0 && local_vf_num == 436 && local_vf_active == 1) port_count[436]++; 
              else if (local_pf_num == 0 && local_vf_num == 437 && local_vf_active == 1) port_count[437]++; 
              else if (local_pf_num == 0 && local_vf_num == 438 && local_vf_active == 1) port_count[438]++; 
              else if (local_pf_num == 0 && local_vf_num == 439 && local_vf_active == 1) port_count[439]++; 
              else if (local_pf_num == 0 && local_vf_num == 440 && local_vf_active == 1) port_count[440]++; 
              else if (local_pf_num == 0 && local_vf_num == 441 && local_vf_active == 1) port_count[441]++; 
              else if (local_pf_num == 0 && local_vf_num == 442 && local_vf_active == 1) port_count[442]++; 
              else if (local_pf_num == 0 && local_vf_num == 443 && local_vf_active == 1) port_count[443]++; 
              else if (local_pf_num == 0 && local_vf_num == 444 && local_vf_active == 1) port_count[444]++; 
              else if (local_pf_num == 0 && local_vf_num == 445 && local_vf_active == 1) port_count[445]++; 
              else if (local_pf_num == 0 && local_vf_num == 446 && local_vf_active == 1) port_count[446]++; 
              else if (local_pf_num == 0 && local_vf_num == 447 && local_vf_active == 1) port_count[447]++; 
              else if (local_pf_num == 0 && local_vf_num == 448 && local_vf_active == 1) port_count[448]++; 
              else if (local_pf_num == 0 && local_vf_num == 449 && local_vf_active == 1) port_count[449]++; 
              else if (local_pf_num == 0 && local_vf_num == 450 && local_vf_active == 1) port_count[450]++; 
              else if (local_pf_num == 0 && local_vf_num == 451 && local_vf_active == 1) port_count[451]++; 
              else if (local_pf_num == 0 && local_vf_num == 452 && local_vf_active == 1) port_count[452]++; 
              else if (local_pf_num == 0 && local_vf_num == 453 && local_vf_active == 1) port_count[453]++; 
              else if (local_pf_num == 0 && local_vf_num == 454 && local_vf_active == 1) port_count[454]++; 
              else if (local_pf_num == 0 && local_vf_num == 455 && local_vf_active == 1) port_count[455]++; 
              else if (local_pf_num == 0 && local_vf_num == 456 && local_vf_active == 1) port_count[456]++; 
              else if (local_pf_num == 0 && local_vf_num == 457 && local_vf_active == 1) port_count[457]++; 
              else if (local_pf_num == 0 && local_vf_num == 458 && local_vf_active == 1) port_count[458]++; 
              else if (local_pf_num == 0 && local_vf_num == 459 && local_vf_active == 1) port_count[459]++; 
              else if (local_pf_num == 0 && local_vf_num == 460 && local_vf_active == 1) port_count[460]++; 
              else if (local_pf_num == 0 && local_vf_num == 461 && local_vf_active == 1) port_count[461]++; 
              else if (local_pf_num == 0 && local_vf_num == 462 && local_vf_active == 1) port_count[462]++; 
              else if (local_pf_num == 0 && local_vf_num == 463 && local_vf_active == 1) port_count[463]++; 
              else if (local_pf_num == 0 && local_vf_num == 464 && local_vf_active == 1) port_count[464]++; 
              else if (local_pf_num == 0 && local_vf_num == 465 && local_vf_active == 1) port_count[465]++; 
              else if (local_pf_num == 0 && local_vf_num == 466 && local_vf_active == 1) port_count[466]++; 
              else if (local_pf_num == 0 && local_vf_num == 467 && local_vf_active == 1) port_count[467]++; 
              else if (local_pf_num == 0 && local_vf_num == 468 && local_vf_active == 1) port_count[468]++; 
              else if (local_pf_num == 0 && local_vf_num == 469 && local_vf_active == 1) port_count[469]++; 
              else if (local_pf_num == 0 && local_vf_num == 470 && local_vf_active == 1) port_count[470]++; 
              else if (local_pf_num == 0 && local_vf_num == 471 && local_vf_active == 1) port_count[471]++; 
              else if (local_pf_num == 0 && local_vf_num == 472 && local_vf_active == 1) port_count[472]++; 
              else if (local_pf_num == 0 && local_vf_num == 473 && local_vf_active == 1) port_count[473]++; 
              else if (local_pf_num == 0 && local_vf_num == 474 && local_vf_active == 1) port_count[474]++; 
              else if (local_pf_num == 0 && local_vf_num == 475 && local_vf_active == 1) port_count[475]++; 
              else if (local_pf_num == 0 && local_vf_num == 476 && local_vf_active == 1) port_count[476]++; 
              else if (local_pf_num == 0 && local_vf_num == 477 && local_vf_active == 1) port_count[477]++; 
              else if (local_pf_num == 0 && local_vf_num == 478 && local_vf_active == 1) port_count[478]++; 
              else if (local_pf_num == 0 && local_vf_num == 479 && local_vf_active == 1) port_count[479]++; 
              else if (local_pf_num == 0 && local_vf_num == 480 && local_vf_active == 1) port_count[480]++; 
              else if (local_pf_num == 0 && local_vf_num == 481 && local_vf_active == 1) port_count[481]++; 
              else if (local_pf_num == 0 && local_vf_num == 482 && local_vf_active == 1) port_count[482]++; 
              else if (local_pf_num == 0 && local_vf_num == 483 && local_vf_active == 1) port_count[483]++; 
              else if (local_pf_num == 0 && local_vf_num == 484 && local_vf_active == 1) port_count[484]++; 
              else if (local_pf_num == 0 && local_vf_num == 485 && local_vf_active == 1) port_count[485]++; 
              else if (local_pf_num == 0 && local_vf_num == 486 && local_vf_active == 1) port_count[486]++; 
              else if (local_pf_num == 0 && local_vf_num == 487 && local_vf_active == 1) port_count[487]++; 
              else if (local_pf_num == 0 && local_vf_num == 488 && local_vf_active == 1) port_count[488]++; 
              else if (local_pf_num == 0 && local_vf_num == 489 && local_vf_active == 1) port_count[489]++; 
              else if (local_pf_num == 0 && local_vf_num == 490 && local_vf_active == 1) port_count[490]++; 
              else if (local_pf_num == 0 && local_vf_num == 491 && local_vf_active == 1) port_count[491]++; 
              else if (local_pf_num == 0 && local_vf_num == 492 && local_vf_active == 1) port_count[492]++; 
              else if (local_pf_num == 0 && local_vf_num == 493 && local_vf_active == 1) port_count[493]++; 
              else if (local_pf_num == 0 && local_vf_num == 494 && local_vf_active == 1) port_count[494]++; 
              else if (local_pf_num == 0 && local_vf_num == 495 && local_vf_active == 1) port_count[495]++; 
              else if (local_pf_num == 0 && local_vf_num == 496 && local_vf_active == 1) port_count[496]++; 
              else if (local_pf_num == 0 && local_vf_num == 497 && local_vf_active == 1) port_count[497]++; 
              else if (local_pf_num == 0 && local_vf_num == 498 && local_vf_active == 1) port_count[498]++; 
              else if (local_pf_num == 0 && local_vf_num == 499 && local_vf_active == 1) port_count[499]++; 
              else if (local_pf_num == 0 && local_vf_num == 500 && local_vf_active == 1) port_count[500]++; 
              else if (local_pf_num == 0 && local_vf_num == 501 && local_vf_active == 1) port_count[501]++; 
              else if (local_pf_num == 0 && local_vf_num == 502 && local_vf_active == 1) port_count[502]++; 
              else if (local_pf_num == 0 && local_vf_num == 503 && local_vf_active == 1) port_count[503]++; 
              else if (local_pf_num == 0 && local_vf_num == 504 && local_vf_active == 1) port_count[504]++; 
              else if (local_pf_num == 0 && local_vf_num == 505 && local_vf_active == 1) port_count[505]++; 
              else if (local_pf_num == 0 && local_vf_num == 506 && local_vf_active == 1) port_count[506]++; 
              else if (local_pf_num == 0 && local_vf_num == 507 && local_vf_active == 1) port_count[507]++; 
              else if (local_pf_num == 0 && local_vf_num == 508 && local_vf_active == 1) port_count[508]++; 
              else if (local_pf_num == 0 && local_vf_num == 509 && local_vf_active == 1) port_count[509]++; 
              else if (local_pf_num == 0 && local_vf_num == 510 && local_vf_active == 1) port_count[510]++; 
              else if (local_pf_num == 0 && local_vf_num == 511 && local_vf_active == 1) port_count[511]++; 
              else if (local_pf_num == 0 && local_vf_num == 512 && local_vf_active == 1) port_count[512]++; 
              else if (local_pf_num == 0 && local_vf_num == 513 && local_vf_active == 1) port_count[513]++; 
              else if (local_pf_num == 0 && local_vf_num == 514 && local_vf_active == 1) port_count[514]++; 
              else if (local_pf_num == 0 && local_vf_num == 515 && local_vf_active == 1) port_count[515]++; 
              else if (local_pf_num == 0 && local_vf_num == 516 && local_vf_active == 1) port_count[516]++; 
              else if (local_pf_num == 0 && local_vf_num == 517 && local_vf_active == 1) port_count[517]++; 
              else if (local_pf_num == 0 && local_vf_num == 518 && local_vf_active == 1) port_count[518]++; 
              else if (local_pf_num == 0 && local_vf_num == 519 && local_vf_active == 1) port_count[519]++; 
              else if (local_pf_num == 0 && local_vf_num == 520 && local_vf_active == 1) port_count[520]++; 
              else if (local_pf_num == 0 && local_vf_num == 521 && local_vf_active == 1) port_count[521]++; 
              else if (local_pf_num == 0 && local_vf_num == 522 && local_vf_active == 1) port_count[522]++; 
              else if (local_pf_num == 0 && local_vf_num == 523 && local_vf_active == 1) port_count[523]++; 
              else if (local_pf_num == 0 && local_vf_num == 524 && local_vf_active == 1) port_count[524]++; 
              else if (local_pf_num == 0 && local_vf_num == 525 && local_vf_active == 1) port_count[525]++; 
              else if (local_pf_num == 0 && local_vf_num == 526 && local_vf_active == 1) port_count[526]++; 
              else if (local_pf_num == 0 && local_vf_num == 527 && local_vf_active == 1) port_count[527]++; 
              else if (local_pf_num == 0 && local_vf_num == 528 && local_vf_active == 1) port_count[528]++; 
              else if (local_pf_num == 0 && local_vf_num == 529 && local_vf_active == 1) port_count[529]++; 
              else if (local_pf_num == 0 && local_vf_num == 530 && local_vf_active == 1) port_count[530]++; 
              else if (local_pf_num == 0 && local_vf_num == 531 && local_vf_active == 1) port_count[531]++; 
              else if (local_pf_num == 0 && local_vf_num == 532 && local_vf_active == 1) port_count[532]++; 
              else if (local_pf_num == 0 && local_vf_num == 533 && local_vf_active == 1) port_count[533]++; 
              else if (local_pf_num == 0 && local_vf_num == 534 && local_vf_active == 1) port_count[534]++; 
              else if (local_pf_num == 0 && local_vf_num == 535 && local_vf_active == 1) port_count[535]++; 
              else if (local_pf_num == 0 && local_vf_num == 536 && local_vf_active == 1) port_count[536]++; 
              else if (local_pf_num == 0 && local_vf_num == 537 && local_vf_active == 1) port_count[537]++; 
              else if (local_pf_num == 0 && local_vf_num == 538 && local_vf_active == 1) port_count[538]++; 
              else if (local_pf_num == 0 && local_vf_num == 539 && local_vf_active == 1) port_count[539]++; 
              else if (local_pf_num == 0 && local_vf_num == 540 && local_vf_active == 1) port_count[540]++; 
              else if (local_pf_num == 0 && local_vf_num == 541 && local_vf_active == 1) port_count[541]++; 
              else if (local_pf_num == 0 && local_vf_num == 542 && local_vf_active == 1) port_count[542]++; 
              else if (local_pf_num == 0 && local_vf_num == 543 && local_vf_active == 1) port_count[543]++; 
              else if (local_pf_num == 0 && local_vf_num == 544 && local_vf_active == 1) port_count[544]++; 
              else if (local_pf_num == 0 && local_vf_num == 545 && local_vf_active == 1) port_count[545]++; 
              else if (local_pf_num == 0 && local_vf_num == 546 && local_vf_active == 1) port_count[546]++; 
              else if (local_pf_num == 0 && local_vf_num == 547 && local_vf_active == 1) port_count[547]++; 
              else if (local_pf_num == 0 && local_vf_num == 548 && local_vf_active == 1) port_count[548]++; 
              else if (local_pf_num == 0 && local_vf_num == 549 && local_vf_active == 1) port_count[549]++; 
              else if (local_pf_num == 0 && local_vf_num == 550 && local_vf_active == 1) port_count[550]++; 
              else if (local_pf_num == 0 && local_vf_num == 551 && local_vf_active == 1) port_count[551]++; 
              else if (local_pf_num == 0 && local_vf_num == 552 && local_vf_active == 1) port_count[552]++; 
              else if (local_pf_num == 0 && local_vf_num == 553 && local_vf_active == 1) port_count[553]++; 
              else if (local_pf_num == 0 && local_vf_num == 554 && local_vf_active == 1) port_count[554]++; 
              else if (local_pf_num == 0 && local_vf_num == 555 && local_vf_active == 1) port_count[555]++; 
              else if (local_pf_num == 0 && local_vf_num == 556 && local_vf_active == 1) port_count[556]++; 
              else if (local_pf_num == 0 && local_vf_num == 557 && local_vf_active == 1) port_count[557]++; 
              else if (local_pf_num == 0 && local_vf_num == 558 && local_vf_active == 1) port_count[558]++; 
              else if (local_pf_num == 0 && local_vf_num == 559 && local_vf_active == 1) port_count[559]++; 
              else if (local_pf_num == 0 && local_vf_num == 560 && local_vf_active == 1) port_count[560]++; 
              else if (local_pf_num == 0 && local_vf_num == 561 && local_vf_active == 1) port_count[561]++; 
              else if (local_pf_num == 0 && local_vf_num == 562 && local_vf_active == 1) port_count[562]++; 
              else if (local_pf_num == 0 && local_vf_num == 563 && local_vf_active == 1) port_count[563]++; 
              else if (local_pf_num == 0 && local_vf_num == 564 && local_vf_active == 1) port_count[564]++; 
              else if (local_pf_num == 0 && local_vf_num == 565 && local_vf_active == 1) port_count[565]++; 
              else if (local_pf_num == 0 && local_vf_num == 566 && local_vf_active == 1) port_count[566]++; 
              else if (local_pf_num == 0 && local_vf_num == 567 && local_vf_active == 1) port_count[567]++; 
              else if (local_pf_num == 0 && local_vf_num == 568 && local_vf_active == 1) port_count[568]++; 
              else if (local_pf_num == 0 && local_vf_num == 569 && local_vf_active == 1) port_count[569]++; 
              else if (local_pf_num == 0 && local_vf_num == 570 && local_vf_active == 1) port_count[570]++; 
              else if (local_pf_num == 0 && local_vf_num == 571 && local_vf_active == 1) port_count[571]++; 
              else if (local_pf_num == 0 && local_vf_num == 572 && local_vf_active == 1) port_count[572]++; 
              else if (local_pf_num == 0 && local_vf_num == 573 && local_vf_active == 1) port_count[573]++; 
              else if (local_pf_num == 0 && local_vf_num == 574 && local_vf_active == 1) port_count[574]++; 
              else if (local_pf_num == 0 && local_vf_num == 575 && local_vf_active == 1) port_count[575]++; 
              else if (local_pf_num == 0 && local_vf_num == 576 && local_vf_active == 1) port_count[576]++; 
              else if (local_pf_num == 0 && local_vf_num == 577 && local_vf_active == 1) port_count[577]++; 
              else if (local_pf_num == 0 && local_vf_num == 578 && local_vf_active == 1) port_count[578]++; 
              else if (local_pf_num == 0 && local_vf_num == 579 && local_vf_active == 1) port_count[579]++; 
              else if (local_pf_num == 0 && local_vf_num == 580 && local_vf_active == 1) port_count[580]++; 
              else if (local_pf_num == 0 && local_vf_num == 581 && local_vf_active == 1) port_count[581]++; 
              else if (local_pf_num == 0 && local_vf_num == 582 && local_vf_active == 1) port_count[582]++; 
              else if (local_pf_num == 0 && local_vf_num == 583 && local_vf_active == 1) port_count[583]++; 
              else if (local_pf_num == 0 && local_vf_num == 584 && local_vf_active == 1) port_count[584]++; 
              else if (local_pf_num == 0 && local_vf_num == 585 && local_vf_active == 1) port_count[585]++; 
              else if (local_pf_num == 0 && local_vf_num == 586 && local_vf_active == 1) port_count[586]++; 
              else if (local_pf_num == 0 && local_vf_num == 587 && local_vf_active == 1) port_count[587]++; 
              else if (local_pf_num == 0 && local_vf_num == 588 && local_vf_active == 1) port_count[588]++; 
              else if (local_pf_num == 0 && local_vf_num == 589 && local_vf_active == 1) port_count[589]++; 
              else if (local_pf_num == 0 && local_vf_num == 590 && local_vf_active == 1) port_count[590]++; 
              else if (local_pf_num == 0 && local_vf_num == 591 && local_vf_active == 1) port_count[591]++; 
              else if (local_pf_num == 0 && local_vf_num == 592 && local_vf_active == 1) port_count[592]++; 
              else if (local_pf_num == 0 && local_vf_num == 593 && local_vf_active == 1) port_count[593]++; 
              else if (local_pf_num == 0 && local_vf_num == 594 && local_vf_active == 1) port_count[594]++; 
              else if (local_pf_num == 0 && local_vf_num == 595 && local_vf_active == 1) port_count[595]++; 
              else if (local_pf_num == 0 && local_vf_num == 596 && local_vf_active == 1) port_count[596]++; 
              else if (local_pf_num == 0 && local_vf_num == 597 && local_vf_active == 1) port_count[597]++; 
              else if (local_pf_num == 0 && local_vf_num == 598 && local_vf_active == 1) port_count[598]++; 
              else if (local_pf_num == 0 && local_vf_num == 599 && local_vf_active == 1) port_count[599]++; 
              else if (local_pf_num == 0 && local_vf_num == 600 && local_vf_active == 1) port_count[600]++; 
              else if (local_pf_num == 0 && local_vf_num == 601 && local_vf_active == 1) port_count[601]++; 
              else if (local_pf_num == 0 && local_vf_num == 602 && local_vf_active == 1) port_count[602]++; 
              else if (local_pf_num == 0 && local_vf_num == 603 && local_vf_active == 1) port_count[603]++; 
              else if (local_pf_num == 0 && local_vf_num == 604 && local_vf_active == 1) port_count[604]++; 
              else if (local_pf_num == 0 && local_vf_num == 605 && local_vf_active == 1) port_count[605]++; 
              else if (local_pf_num == 0 && local_vf_num == 606 && local_vf_active == 1) port_count[606]++; 
              else if (local_pf_num == 0 && local_vf_num == 607 && local_vf_active == 1) port_count[607]++; 
              else if (local_pf_num == 0 && local_vf_num == 608 && local_vf_active == 1) port_count[608]++; 
              else if (local_pf_num == 0 && local_vf_num == 609 && local_vf_active == 1) port_count[609]++; 
              else if (local_pf_num == 0 && local_vf_num == 610 && local_vf_active == 1) port_count[610]++; 
              else if (local_pf_num == 0 && local_vf_num == 611 && local_vf_active == 1) port_count[611]++; 
              else if (local_pf_num == 0 && local_vf_num == 612 && local_vf_active == 1) port_count[612]++; 
              else if (local_pf_num == 0 && local_vf_num == 613 && local_vf_active == 1) port_count[613]++; 
              else if (local_pf_num == 0 && local_vf_num == 614 && local_vf_active == 1) port_count[614]++; 
              else if (local_pf_num == 0 && local_vf_num == 615 && local_vf_active == 1) port_count[615]++; 
              else if (local_pf_num == 0 && local_vf_num == 616 && local_vf_active == 1) port_count[616]++; 
              else if (local_pf_num == 0 && local_vf_num == 617 && local_vf_active == 1) port_count[617]++; 
              else if (local_pf_num == 0 && local_vf_num == 618 && local_vf_active == 1) port_count[618]++; 
              else if (local_pf_num == 0 && local_vf_num == 619 && local_vf_active == 1) port_count[619]++; 
              else if (local_pf_num == 0 && local_vf_num == 620 && local_vf_active == 1) port_count[620]++; 
              else if (local_pf_num == 0 && local_vf_num == 621 && local_vf_active == 1) port_count[621]++; 
              else if (local_pf_num == 0 && local_vf_num == 622 && local_vf_active == 1) port_count[622]++; 
              else if (local_pf_num == 0 && local_vf_num == 623 && local_vf_active == 1) port_count[623]++; 
              else if (local_pf_num == 0 && local_vf_num == 624 && local_vf_active == 1) port_count[624]++; 
              else if (local_pf_num == 0 && local_vf_num == 625 && local_vf_active == 1) port_count[625]++; 
              else if (local_pf_num == 0 && local_vf_num == 626 && local_vf_active == 1) port_count[626]++; 
              else if (local_pf_num == 0 && local_vf_num == 627 && local_vf_active == 1) port_count[627]++; 
              else if (local_pf_num == 0 && local_vf_num == 628 && local_vf_active == 1) port_count[628]++; 
              else if (local_pf_num == 0 && local_vf_num == 629 && local_vf_active == 1) port_count[629]++; 
              else if (local_pf_num == 0 && local_vf_num == 630 && local_vf_active == 1) port_count[630]++; 
              else if (local_pf_num == 0 && local_vf_num == 631 && local_vf_active == 1) port_count[631]++; 
              else if (local_pf_num == 0 && local_vf_num == 632 && local_vf_active == 1) port_count[632]++; 
              else if (local_pf_num == 0 && local_vf_num == 633 && local_vf_active == 1) port_count[633]++; 
              else if (local_pf_num == 0 && local_vf_num == 634 && local_vf_active == 1) port_count[634]++; 
              else if (local_pf_num == 0 && local_vf_num == 635 && local_vf_active == 1) port_count[635]++; 
              else if (local_pf_num == 0 && local_vf_num == 636 && local_vf_active == 1) port_count[636]++; 
              else if (local_pf_num == 0 && local_vf_num == 637 && local_vf_active == 1) port_count[637]++; 
              else if (local_pf_num == 0 && local_vf_num == 638 && local_vf_active == 1) port_count[638]++; 
              else if (local_pf_num == 0 && local_vf_num == 639 && local_vf_active == 1) port_count[639]++; 
              else if (local_pf_num == 0 && local_vf_num == 640 && local_vf_active == 1) port_count[640]++; 
              else if (local_pf_num == 0 && local_vf_num == 641 && local_vf_active == 1) port_count[641]++; 
              else if (local_pf_num == 0 && local_vf_num == 642 && local_vf_active == 1) port_count[642]++; 
              else if (local_pf_num == 0 && local_vf_num == 643 && local_vf_active == 1) port_count[643]++; 
              else if (local_pf_num == 0 && local_vf_num == 644 && local_vf_active == 1) port_count[644]++; 
              else if (local_pf_num == 0 && local_vf_num == 645 && local_vf_active == 1) port_count[645]++; 
              else if (local_pf_num == 0 && local_vf_num == 646 && local_vf_active == 1) port_count[646]++; 
              else if (local_pf_num == 0 && local_vf_num == 647 && local_vf_active == 1) port_count[647]++; 
              else if (local_pf_num == 0 && local_vf_num == 648 && local_vf_active == 1) port_count[648]++; 
              else if (local_pf_num == 0 && local_vf_num == 649 && local_vf_active == 1) port_count[649]++; 
              else if (local_pf_num == 0 && local_vf_num == 650 && local_vf_active == 1) port_count[650]++; 
              else if (local_pf_num == 0 && local_vf_num == 651 && local_vf_active == 1) port_count[651]++; 
              else if (local_pf_num == 0 && local_vf_num == 652 && local_vf_active == 1) port_count[652]++; 
              else if (local_pf_num == 0 && local_vf_num == 653 && local_vf_active == 1) port_count[653]++; 
              else if (local_pf_num == 0 && local_vf_num == 654 && local_vf_active == 1) port_count[654]++; 
              else if (local_pf_num == 0 && local_vf_num == 655 && local_vf_active == 1) port_count[655]++; 
              else if (local_pf_num == 0 && local_vf_num == 656 && local_vf_active == 1) port_count[656]++; 
              else if (local_pf_num == 0 && local_vf_num == 657 && local_vf_active == 1) port_count[657]++; 
              else if (local_pf_num == 0 && local_vf_num == 658 && local_vf_active == 1) port_count[658]++; 
              else if (local_pf_num == 0 && local_vf_num == 659 && local_vf_active == 1) port_count[659]++; 
              else if (local_pf_num == 0 && local_vf_num == 660 && local_vf_active == 1) port_count[660]++; 
              else if (local_pf_num == 0 && local_vf_num == 661 && local_vf_active == 1) port_count[661]++; 
              else if (local_pf_num == 0 && local_vf_num == 662 && local_vf_active == 1) port_count[662]++; 
              else if (local_pf_num == 0 && local_vf_num == 663 && local_vf_active == 1) port_count[663]++; 
              else if (local_pf_num == 0 && local_vf_num == 664 && local_vf_active == 1) port_count[664]++; 
              else if (local_pf_num == 0 && local_vf_num == 665 && local_vf_active == 1) port_count[665]++; 
              else if (local_pf_num == 0 && local_vf_num == 666 && local_vf_active == 1) port_count[666]++; 
              else if (local_pf_num == 0 && local_vf_num == 667 && local_vf_active == 1) port_count[667]++; 
              else if (local_pf_num == 0 && local_vf_num == 668 && local_vf_active == 1) port_count[668]++; 
              else if (local_pf_num == 0 && local_vf_num == 669 && local_vf_active == 1) port_count[669]++; 
              else if (local_pf_num == 0 && local_vf_num == 670 && local_vf_active == 1) port_count[670]++; 
              else if (local_pf_num == 0 && local_vf_num == 671 && local_vf_active == 1) port_count[671]++; 
              else if (local_pf_num == 0 && local_vf_num == 672 && local_vf_active == 1) port_count[672]++; 
              else if (local_pf_num == 0 && local_vf_num == 673 && local_vf_active == 1) port_count[673]++; 
              else if (local_pf_num == 0 && local_vf_num == 674 && local_vf_active == 1) port_count[674]++; 
              else if (local_pf_num == 0 && local_vf_num == 675 && local_vf_active == 1) port_count[675]++; 
              else if (local_pf_num == 0 && local_vf_num == 676 && local_vf_active == 1) port_count[676]++; 
              else if (local_pf_num == 0 && local_vf_num == 677 && local_vf_active == 1) port_count[677]++; 
              else if (local_pf_num == 0 && local_vf_num == 678 && local_vf_active == 1) port_count[678]++; 
              else if (local_pf_num == 0 && local_vf_num == 679 && local_vf_active == 1) port_count[679]++; 
              else if (local_pf_num == 0 && local_vf_num == 680 && local_vf_active == 1) port_count[680]++; 
              else if (local_pf_num == 0 && local_vf_num == 681 && local_vf_active == 1) port_count[681]++; 
              else if (local_pf_num == 0 && local_vf_num == 682 && local_vf_active == 1) port_count[682]++; 
              else if (local_pf_num == 0 && local_vf_num == 683 && local_vf_active == 1) port_count[683]++; 
              else if (local_pf_num == 0 && local_vf_num == 684 && local_vf_active == 1) port_count[684]++; 
              else if (local_pf_num == 0 && local_vf_num == 685 && local_vf_active == 1) port_count[685]++; 
              else if (local_pf_num == 0 && local_vf_num == 686 && local_vf_active == 1) port_count[686]++; 
              else if (local_pf_num == 0 && local_vf_num == 687 && local_vf_active == 1) port_count[687]++; 
              else if (local_pf_num == 0 && local_vf_num == 688 && local_vf_active == 1) port_count[688]++; 
              else if (local_pf_num == 0 && local_vf_num == 689 && local_vf_active == 1) port_count[689]++; 
              else if (local_pf_num == 0 && local_vf_num == 690 && local_vf_active == 1) port_count[690]++; 
              else if (local_pf_num == 0 && local_vf_num == 691 && local_vf_active == 1) port_count[691]++; 
              else if (local_pf_num == 0 && local_vf_num == 692 && local_vf_active == 1) port_count[692]++; 
              else if (local_pf_num == 0 && local_vf_num == 693 && local_vf_active == 1) port_count[693]++; 
              else if (local_pf_num == 0 && local_vf_num == 694 && local_vf_active == 1) port_count[694]++; 
              else if (local_pf_num == 0 && local_vf_num == 695 && local_vf_active == 1) port_count[695]++; 
              else if (local_pf_num == 0 && local_vf_num == 696 && local_vf_active == 1) port_count[696]++; 
              else if (local_pf_num == 0 && local_vf_num == 697 && local_vf_active == 1) port_count[697]++; 
              else if (local_pf_num == 0 && local_vf_num == 698 && local_vf_active == 1) port_count[698]++; 
              else if (local_pf_num == 0 && local_vf_num == 699 && local_vf_active == 1) port_count[699]++; 
              else if (local_pf_num == 0 && local_vf_num == 700 && local_vf_active == 1) port_count[700]++; 
              else if (local_pf_num == 0 && local_vf_num == 701 && local_vf_active == 1) port_count[701]++; 
              else if (local_pf_num == 0 && local_vf_num == 702 && local_vf_active == 1) port_count[702]++; 
              else if (local_pf_num == 0 && local_vf_num == 703 && local_vf_active == 1) port_count[703]++; 
              else if (local_pf_num == 0 && local_vf_num == 704 && local_vf_active == 1) port_count[704]++; 
              else if (local_pf_num == 0 && local_vf_num == 705 && local_vf_active == 1) port_count[705]++; 
              else if (local_pf_num == 0 && local_vf_num == 706 && local_vf_active == 1) port_count[706]++; 
              else if (local_pf_num == 0 && local_vf_num == 707 && local_vf_active == 1) port_count[707]++; 
              else if (local_pf_num == 0 && local_vf_num == 708 && local_vf_active == 1) port_count[708]++; 
              else if (local_pf_num == 0 && local_vf_num == 709 && local_vf_active == 1) port_count[709]++; 
              else if (local_pf_num == 0 && local_vf_num == 710 && local_vf_active == 1) port_count[710]++; 
              else if (local_pf_num == 0 && local_vf_num == 711 && local_vf_active == 1) port_count[711]++; 
              else if (local_pf_num == 0 && local_vf_num == 712 && local_vf_active == 1) port_count[712]++; 
              else if (local_pf_num == 0 && local_vf_num == 713 && local_vf_active == 1) port_count[713]++; 
              else if (local_pf_num == 0 && local_vf_num == 714 && local_vf_active == 1) port_count[714]++; 
              else if (local_pf_num == 0 && local_vf_num == 715 && local_vf_active == 1) port_count[715]++; 
              else if (local_pf_num == 0 && local_vf_num == 716 && local_vf_active == 1) port_count[716]++; 
              else if (local_pf_num == 0 && local_vf_num == 717 && local_vf_active == 1) port_count[717]++; 
              else if (local_pf_num == 0 && local_vf_num == 718 && local_vf_active == 1) port_count[718]++; 
              else if (local_pf_num == 0 && local_vf_num == 719 && local_vf_active == 1) port_count[719]++; 
              else if (local_pf_num == 0 && local_vf_num == 720 && local_vf_active == 1) port_count[720]++; 
              else if (local_pf_num == 0 && local_vf_num == 721 && local_vf_active == 1) port_count[721]++; 
              else if (local_pf_num == 0 && local_vf_num == 722 && local_vf_active == 1) port_count[722]++; 
              else if (local_pf_num == 0 && local_vf_num == 723 && local_vf_active == 1) port_count[723]++; 
              else if (local_pf_num == 0 && local_vf_num == 724 && local_vf_active == 1) port_count[724]++; 
              else if (local_pf_num == 0 && local_vf_num == 725 && local_vf_active == 1) port_count[725]++; 
              else if (local_pf_num == 0 && local_vf_num == 726 && local_vf_active == 1) port_count[726]++; 
              else if (local_pf_num == 0 && local_vf_num == 727 && local_vf_active == 1) port_count[727]++; 
              else if (local_pf_num == 0 && local_vf_num == 728 && local_vf_active == 1) port_count[728]++; 
              else if (local_pf_num == 0 && local_vf_num == 729 && local_vf_active == 1) port_count[729]++; 
              else if (local_pf_num == 0 && local_vf_num == 730 && local_vf_active == 1) port_count[730]++; 
              else if (local_pf_num == 0 && local_vf_num == 731 && local_vf_active == 1) port_count[731]++; 
              else if (local_pf_num == 0 && local_vf_num == 732 && local_vf_active == 1) port_count[732]++; 
              else if (local_pf_num == 0 && local_vf_num == 733 && local_vf_active == 1) port_count[733]++; 
              else if (local_pf_num == 0 && local_vf_num == 734 && local_vf_active == 1) port_count[734]++; 
              else if (local_pf_num == 0 && local_vf_num == 735 && local_vf_active == 1) port_count[735]++; 
              else if (local_pf_num == 0 && local_vf_num == 736 && local_vf_active == 1) port_count[736]++; 
              else if (local_pf_num == 0 && local_vf_num == 737 && local_vf_active == 1) port_count[737]++; 
              else if (local_pf_num == 0 && local_vf_num == 738 && local_vf_active == 1) port_count[738]++; 
              else if (local_pf_num == 0 && local_vf_num == 739 && local_vf_active == 1) port_count[739]++; 
              else if (local_pf_num == 0 && local_vf_num == 740 && local_vf_active == 1) port_count[740]++; 
              else if (local_pf_num == 0 && local_vf_num == 741 && local_vf_active == 1) port_count[741]++; 
              else if (local_pf_num == 0 && local_vf_num == 742 && local_vf_active == 1) port_count[742]++; 
              else if (local_pf_num == 0 && local_vf_num == 743 && local_vf_active == 1) port_count[743]++; 
              else if (local_pf_num == 0 && local_vf_num == 744 && local_vf_active == 1) port_count[744]++; 
              else if (local_pf_num == 0 && local_vf_num == 745 && local_vf_active == 1) port_count[745]++; 
              else if (local_pf_num == 0 && local_vf_num == 746 && local_vf_active == 1) port_count[746]++; 
              else if (local_pf_num == 0 && local_vf_num == 747 && local_vf_active == 1) port_count[747]++; 
              else if (local_pf_num == 0 && local_vf_num == 748 && local_vf_active == 1) port_count[748]++; 
              else if (local_pf_num == 0 && local_vf_num == 749 && local_vf_active == 1) port_count[749]++; 
              else if (local_pf_num == 0 && local_vf_num == 750 && local_vf_active == 1) port_count[750]++; 
              else if (local_pf_num == 0 && local_vf_num == 751 && local_vf_active == 1) port_count[751]++; 
              else if (local_pf_num == 0 && local_vf_num == 752 && local_vf_active == 1) port_count[752]++; 
              else if (local_pf_num == 0 && local_vf_num == 753 && local_vf_active == 1) port_count[753]++; 
              else if (local_pf_num == 0 && local_vf_num == 754 && local_vf_active == 1) port_count[754]++; 
              else if (local_pf_num == 0 && local_vf_num == 755 && local_vf_active == 1) port_count[755]++; 
              else if (local_pf_num == 0 && local_vf_num == 756 && local_vf_active == 1) port_count[756]++; 
              else if (local_pf_num == 0 && local_vf_num == 757 && local_vf_active == 1) port_count[757]++; 
              else if (local_pf_num == 0 && local_vf_num == 758 && local_vf_active == 1) port_count[758]++; 
              else if (local_pf_num == 0 && local_vf_num == 759 && local_vf_active == 1) port_count[759]++; 
              else if (local_pf_num == 0 && local_vf_num == 760 && local_vf_active == 1) port_count[760]++; 
              else if (local_pf_num == 0 && local_vf_num == 761 && local_vf_active == 1) port_count[761]++; 
              else if (local_pf_num == 0 && local_vf_num == 762 && local_vf_active == 1) port_count[762]++; 
              else if (local_pf_num == 0 && local_vf_num == 763 && local_vf_active == 1) port_count[763]++; 
              else if (local_pf_num == 0 && local_vf_num == 764 && local_vf_active == 1) port_count[764]++; 
              else if (local_pf_num == 0 && local_vf_num == 765 && local_vf_active == 1) port_count[765]++; 
              else if (local_pf_num == 0 && local_vf_num == 766 && local_vf_active == 1) port_count[766]++; 
              else if (local_pf_num == 0 && local_vf_num == 767 && local_vf_active == 1) port_count[767]++; 
              else if (local_pf_num == 0 && local_vf_num == 768 && local_vf_active == 1) port_count[768]++; 
              else if (local_pf_num == 0 && local_vf_num == 769 && local_vf_active == 1) port_count[769]++; 
              else if (local_pf_num == 0 && local_vf_num == 770 && local_vf_active == 1) port_count[770]++; 
              else if (local_pf_num == 0 && local_vf_num == 771 && local_vf_active == 1) port_count[771]++; 
              else if (local_pf_num == 0 && local_vf_num == 772 && local_vf_active == 1) port_count[772]++; 
              else if (local_pf_num == 0 && local_vf_num == 773 && local_vf_active == 1) port_count[773]++; 
              else if (local_pf_num == 0 && local_vf_num == 774 && local_vf_active == 1) port_count[774]++; 
              else if (local_pf_num == 0 && local_vf_num == 775 && local_vf_active == 1) port_count[775]++; 
              else if (local_pf_num == 0 && local_vf_num == 776 && local_vf_active == 1) port_count[776]++; 
              else if (local_pf_num == 0 && local_vf_num == 777 && local_vf_active == 1) port_count[777]++; 
              else if (local_pf_num == 0 && local_vf_num == 778 && local_vf_active == 1) port_count[778]++; 
              else if (local_pf_num == 0 && local_vf_num == 779 && local_vf_active == 1) port_count[779]++; 
              else if (local_pf_num == 0 && local_vf_num == 780 && local_vf_active == 1) port_count[780]++; 
              else if (local_pf_num == 0 && local_vf_num == 781 && local_vf_active == 1) port_count[781]++; 
              else if (local_pf_num == 0 && local_vf_num == 782 && local_vf_active == 1) port_count[782]++; 
              else if (local_pf_num == 0 && local_vf_num == 783 && local_vf_active == 1) port_count[783]++; 
              else if (local_pf_num == 0 && local_vf_num == 784 && local_vf_active == 1) port_count[784]++; 
              else if (local_pf_num == 0 && local_vf_num == 785 && local_vf_active == 1) port_count[785]++; 
              else if (local_pf_num == 0 && local_vf_num == 786 && local_vf_active == 1) port_count[786]++; 
              else if (local_pf_num == 0 && local_vf_num == 787 && local_vf_active == 1) port_count[787]++; 
              else if (local_pf_num == 0 && local_vf_num == 788 && local_vf_active == 1) port_count[788]++; 
              else if (local_pf_num == 0 && local_vf_num == 789 && local_vf_active == 1) port_count[789]++; 
              else if (local_pf_num == 0 && local_vf_num == 790 && local_vf_active == 1) port_count[790]++; 
              else if (local_pf_num == 0 && local_vf_num == 791 && local_vf_active == 1) port_count[791]++; 
              else if (local_pf_num == 0 && local_vf_num == 792 && local_vf_active == 1) port_count[792]++; 
              else if (local_pf_num == 0 && local_vf_num == 793 && local_vf_active == 1) port_count[793]++; 
              else if (local_pf_num == 0 && local_vf_num == 794 && local_vf_active == 1) port_count[794]++; 
              else if (local_pf_num == 0 && local_vf_num == 795 && local_vf_active == 1) port_count[795]++; 
              else if (local_pf_num == 0 && local_vf_num == 796 && local_vf_active == 1) port_count[796]++; 
              else if (local_pf_num == 0 && local_vf_num == 797 && local_vf_active == 1) port_count[797]++; 
              else if (local_pf_num == 0 && local_vf_num == 798 && local_vf_active == 1) port_count[798]++; 
              else if (local_pf_num == 0 && local_vf_num == 799 && local_vf_active == 1) port_count[799]++; 
              else if (local_pf_num == 0 && local_vf_num == 800 && local_vf_active == 1) port_count[800]++; 
              else if (local_pf_num == 0 && local_vf_num == 801 && local_vf_active == 1) port_count[801]++; 
              else if (local_pf_num == 0 && local_vf_num == 802 && local_vf_active == 1) port_count[802]++; 
              else if (local_pf_num == 0 && local_vf_num == 803 && local_vf_active == 1) port_count[803]++; 
              else if (local_pf_num == 0 && local_vf_num == 804 && local_vf_active == 1) port_count[804]++; 
              else if (local_pf_num == 0 && local_vf_num == 805 && local_vf_active == 1) port_count[805]++; 
              else if (local_pf_num == 0 && local_vf_num == 806 && local_vf_active == 1) port_count[806]++; 
              else if (local_pf_num == 0 && local_vf_num == 807 && local_vf_active == 1) port_count[807]++; 
              else if (local_pf_num == 0 && local_vf_num == 808 && local_vf_active == 1) port_count[808]++; 
              else if (local_pf_num == 0 && local_vf_num == 809 && local_vf_active == 1) port_count[809]++; 
              else if (local_pf_num == 0 && local_vf_num == 810 && local_vf_active == 1) port_count[810]++; 
              else if (local_pf_num == 0 && local_vf_num == 811 && local_vf_active == 1) port_count[811]++; 
              else if (local_pf_num == 0 && local_vf_num == 812 && local_vf_active == 1) port_count[812]++; 
              else if (local_pf_num == 0 && local_vf_num == 813 && local_vf_active == 1) port_count[813]++; 
              else if (local_pf_num == 0 && local_vf_num == 814 && local_vf_active == 1) port_count[814]++; 
              else if (local_pf_num == 0 && local_vf_num == 815 && local_vf_active == 1) port_count[815]++; 
              else if (local_pf_num == 0 && local_vf_num == 816 && local_vf_active == 1) port_count[816]++; 
              else if (local_pf_num == 0 && local_vf_num == 817 && local_vf_active == 1) port_count[817]++; 
              else if (local_pf_num == 0 && local_vf_num == 818 && local_vf_active == 1) port_count[818]++; 
              else if (local_pf_num == 0 && local_vf_num == 819 && local_vf_active == 1) port_count[819]++; 
              else if (local_pf_num == 0 && local_vf_num == 820 && local_vf_active == 1) port_count[820]++; 
              else if (local_pf_num == 0 && local_vf_num == 821 && local_vf_active == 1) port_count[821]++; 
              else if (local_pf_num == 0 && local_vf_num == 822 && local_vf_active == 1) port_count[822]++; 
              else if (local_pf_num == 0 && local_vf_num == 823 && local_vf_active == 1) port_count[823]++; 
              else if (local_pf_num == 0 && local_vf_num == 824 && local_vf_active == 1) port_count[824]++; 
              else if (local_pf_num == 0 && local_vf_num == 825 && local_vf_active == 1) port_count[825]++; 
              else if (local_pf_num == 0 && local_vf_num == 826 && local_vf_active == 1) port_count[826]++; 
              else if (local_pf_num == 0 && local_vf_num == 827 && local_vf_active == 1) port_count[827]++; 
              else if (local_pf_num == 0 && local_vf_num == 828 && local_vf_active == 1) port_count[828]++; 
              else if (local_pf_num == 0 && local_vf_num == 829 && local_vf_active == 1) port_count[829]++; 
              else if (local_pf_num == 0 && local_vf_num == 830 && local_vf_active == 1) port_count[830]++; 
              else if (local_pf_num == 0 && local_vf_num == 831 && local_vf_active == 1) port_count[831]++; 
              else if (local_pf_num == 0 && local_vf_num == 832 && local_vf_active == 1) port_count[832]++; 
              else if (local_pf_num == 0 && local_vf_num == 833 && local_vf_active == 1) port_count[833]++; 
              else if (local_pf_num == 0 && local_vf_num == 834 && local_vf_active == 1) port_count[834]++; 
              else if (local_pf_num == 0 && local_vf_num == 835 && local_vf_active == 1) port_count[835]++; 
              else if (local_pf_num == 0 && local_vf_num == 836 && local_vf_active == 1) port_count[836]++; 
              else if (local_pf_num == 0 && local_vf_num == 837 && local_vf_active == 1) port_count[837]++; 
              else if (local_pf_num == 0 && local_vf_num == 838 && local_vf_active == 1) port_count[838]++; 
              else if (local_pf_num == 0 && local_vf_num == 839 && local_vf_active == 1) port_count[839]++; 
              else if (local_pf_num == 0 && local_vf_num == 840 && local_vf_active == 1) port_count[840]++; 
              else if (local_pf_num == 0 && local_vf_num == 841 && local_vf_active == 1) port_count[841]++; 
              else if (local_pf_num == 0 && local_vf_num == 842 && local_vf_active == 1) port_count[842]++; 
              else if (local_pf_num == 0 && local_vf_num == 843 && local_vf_active == 1) port_count[843]++; 
              else if (local_pf_num == 0 && local_vf_num == 844 && local_vf_active == 1) port_count[844]++; 
              else if (local_pf_num == 0 && local_vf_num == 845 && local_vf_active == 1) port_count[845]++; 
              else if (local_pf_num == 0 && local_vf_num == 846 && local_vf_active == 1) port_count[846]++; 
              else if (local_pf_num == 0 && local_vf_num == 847 && local_vf_active == 1) port_count[847]++; 
              else if (local_pf_num == 0 && local_vf_num == 848 && local_vf_active == 1) port_count[848]++; 
              else if (local_pf_num == 0 && local_vf_num == 849 && local_vf_active == 1) port_count[849]++; 
              else if (local_pf_num == 0 && local_vf_num == 850 && local_vf_active == 1) port_count[850]++; 
              else if (local_pf_num == 0 && local_vf_num == 851 && local_vf_active == 1) port_count[851]++; 
              else if (local_pf_num == 0 && local_vf_num == 852 && local_vf_active == 1) port_count[852]++; 
              else if (local_pf_num == 0 && local_vf_num == 853 && local_vf_active == 1) port_count[853]++; 
              else if (local_pf_num == 0 && local_vf_num == 854 && local_vf_active == 1) port_count[854]++; 
              else if (local_pf_num == 0 && local_vf_num == 855 && local_vf_active == 1) port_count[855]++; 
              else if (local_pf_num == 0 && local_vf_num == 856 && local_vf_active == 1) port_count[856]++; 
              else if (local_pf_num == 0 && local_vf_num == 857 && local_vf_active == 1) port_count[857]++; 
              else if (local_pf_num == 0 && local_vf_num == 858 && local_vf_active == 1) port_count[858]++; 
              else if (local_pf_num == 0 && local_vf_num == 859 && local_vf_active == 1) port_count[859]++; 
              else if (local_pf_num == 0 && local_vf_num == 860 && local_vf_active == 1) port_count[860]++; 
              else if (local_pf_num == 0 && local_vf_num == 861 && local_vf_active == 1) port_count[861]++; 
              else if (local_pf_num == 0 && local_vf_num == 862 && local_vf_active == 1) port_count[862]++; 
              else if (local_pf_num == 0 && local_vf_num == 863 && local_vf_active == 1) port_count[863]++; 
              else if (local_pf_num == 0 && local_vf_num == 864 && local_vf_active == 1) port_count[864]++; 
              else if (local_pf_num == 0 && local_vf_num == 865 && local_vf_active == 1) port_count[865]++; 
              else if (local_pf_num == 0 && local_vf_num == 866 && local_vf_active == 1) port_count[866]++; 
              else if (local_pf_num == 0 && local_vf_num == 867 && local_vf_active == 1) port_count[867]++; 
              else if (local_pf_num == 0 && local_vf_num == 868 && local_vf_active == 1) port_count[868]++; 
              else if (local_pf_num == 0 && local_vf_num == 869 && local_vf_active == 1) port_count[869]++; 
              else if (local_pf_num == 0 && local_vf_num == 870 && local_vf_active == 1) port_count[870]++; 
              else if (local_pf_num == 0 && local_vf_num == 871 && local_vf_active == 1) port_count[871]++; 
              else if (local_pf_num == 0 && local_vf_num == 872 && local_vf_active == 1) port_count[872]++; 
              else if (local_pf_num == 0 && local_vf_num == 873 && local_vf_active == 1) port_count[873]++; 
              else if (local_pf_num == 0 && local_vf_num == 874 && local_vf_active == 1) port_count[874]++; 
              else if (local_pf_num == 0 && local_vf_num == 875 && local_vf_active == 1) port_count[875]++; 
              else if (local_pf_num == 0 && local_vf_num == 876 && local_vf_active == 1) port_count[876]++; 
              else if (local_pf_num == 0 && local_vf_num == 877 && local_vf_active == 1) port_count[877]++; 
              else if (local_pf_num == 0 && local_vf_num == 878 && local_vf_active == 1) port_count[878]++; 
              else if (local_pf_num == 0 && local_vf_num == 879 && local_vf_active == 1) port_count[879]++; 
              else if (local_pf_num == 0 && local_vf_num == 880 && local_vf_active == 1) port_count[880]++; 
              else if (local_pf_num == 0 && local_vf_num == 881 && local_vf_active == 1) port_count[881]++; 
              else if (local_pf_num == 0 && local_vf_num == 882 && local_vf_active == 1) port_count[882]++; 
              else if (local_pf_num == 0 && local_vf_num == 883 && local_vf_active == 1) port_count[883]++; 
              else if (local_pf_num == 0 && local_vf_num == 884 && local_vf_active == 1) port_count[884]++; 
              else if (local_pf_num == 0 && local_vf_num == 885 && local_vf_active == 1) port_count[885]++; 
              else if (local_pf_num == 0 && local_vf_num == 886 && local_vf_active == 1) port_count[886]++; 
              else if (local_pf_num == 0 && local_vf_num == 887 && local_vf_active == 1) port_count[887]++; 
              else if (local_pf_num == 0 && local_vf_num == 888 && local_vf_active == 1) port_count[888]++; 
              else if (local_pf_num == 0 && local_vf_num == 889 && local_vf_active == 1) port_count[889]++; 
              else if (local_pf_num == 0 && local_vf_num == 890 && local_vf_active == 1) port_count[890]++; 
              else if (local_pf_num == 0 && local_vf_num == 891 && local_vf_active == 1) port_count[891]++; 
              else if (local_pf_num == 0 && local_vf_num == 892 && local_vf_active == 1) port_count[892]++; 
              else if (local_pf_num == 0 && local_vf_num == 893 && local_vf_active == 1) port_count[893]++; 
              else if (local_pf_num == 0 && local_vf_num == 894 && local_vf_active == 1) port_count[894]++; 
              else if (local_pf_num == 0 && local_vf_num == 895 && local_vf_active == 1) port_count[895]++; 
              else if (local_pf_num == 0 && local_vf_num == 896 && local_vf_active == 1) port_count[896]++; 
              else if (local_pf_num == 0 && local_vf_num == 897 && local_vf_active == 1) port_count[897]++; 
              else if (local_pf_num == 0 && local_vf_num == 898 && local_vf_active == 1) port_count[898]++; 
              else if (local_pf_num == 0 && local_vf_num == 899 && local_vf_active == 1) port_count[899]++; 
              else if (local_pf_num == 0 && local_vf_num == 900 && local_vf_active == 1) port_count[900]++; 
              else if (local_pf_num == 0 && local_vf_num == 901 && local_vf_active == 1) port_count[901]++; 
              else if (local_pf_num == 0 && local_vf_num == 902 && local_vf_active == 1) port_count[902]++; 
              else if (local_pf_num == 0 && local_vf_num == 903 && local_vf_active == 1) port_count[903]++; 
              else if (local_pf_num == 0 && local_vf_num == 904 && local_vf_active == 1) port_count[904]++; 
              else if (local_pf_num == 0 && local_vf_num == 905 && local_vf_active == 1) port_count[905]++; 
              else if (local_pf_num == 0 && local_vf_num == 906 && local_vf_active == 1) port_count[906]++; 
              else if (local_pf_num == 0 && local_vf_num == 907 && local_vf_active == 1) port_count[907]++; 
              else if (local_pf_num == 0 && local_vf_num == 908 && local_vf_active == 1) port_count[908]++; 
              else if (local_pf_num == 0 && local_vf_num == 909 && local_vf_active == 1) port_count[909]++; 
              else if (local_pf_num == 0 && local_vf_num == 910 && local_vf_active == 1) port_count[910]++; 
              else if (local_pf_num == 0 && local_vf_num == 911 && local_vf_active == 1) port_count[911]++; 
              else if (local_pf_num == 0 && local_vf_num == 912 && local_vf_active == 1) port_count[912]++; 
              else if (local_pf_num == 0 && local_vf_num == 913 && local_vf_active == 1) port_count[913]++; 
              else if (local_pf_num == 0 && local_vf_num == 914 && local_vf_active == 1) port_count[914]++; 
              else if (local_pf_num == 0 && local_vf_num == 915 && local_vf_active == 1) port_count[915]++; 
              else if (local_pf_num == 0 && local_vf_num == 916 && local_vf_active == 1) port_count[916]++; 
              else if (local_pf_num == 0 && local_vf_num == 917 && local_vf_active == 1) port_count[917]++; 
              else if (local_pf_num == 0 && local_vf_num == 918 && local_vf_active == 1) port_count[918]++; 
              else if (local_pf_num == 0 && local_vf_num == 919 && local_vf_active == 1) port_count[919]++; 
              else if (local_pf_num == 0 && local_vf_num == 920 && local_vf_active == 1) port_count[920]++; 
              else if (local_pf_num == 0 && local_vf_num == 921 && local_vf_active == 1) port_count[921]++; 
              else if (local_pf_num == 0 && local_vf_num == 922 && local_vf_active == 1) port_count[922]++; 
              else if (local_pf_num == 0 && local_vf_num == 923 && local_vf_active == 1) port_count[923]++; 
              else if (local_pf_num == 0 && local_vf_num == 924 && local_vf_active == 1) port_count[924]++; 
              else if (local_pf_num == 0 && local_vf_num == 925 && local_vf_active == 1) port_count[925]++; 
              else if (local_pf_num == 0 && local_vf_num == 926 && local_vf_active == 1) port_count[926]++; 
              else if (local_pf_num == 0 && local_vf_num == 927 && local_vf_active == 1) port_count[927]++; 
              else if (local_pf_num == 0 && local_vf_num == 928 && local_vf_active == 1) port_count[928]++; 
              else if (local_pf_num == 0 && local_vf_num == 929 && local_vf_active == 1) port_count[929]++; 
              else if (local_pf_num == 0 && local_vf_num == 930 && local_vf_active == 1) port_count[930]++; 
              else if (local_pf_num == 0 && local_vf_num == 931 && local_vf_active == 1) port_count[931]++; 
              else if (local_pf_num == 0 && local_vf_num == 932 && local_vf_active == 1) port_count[932]++; 
              else if (local_pf_num == 0 && local_vf_num == 933 && local_vf_active == 1) port_count[933]++; 
              else if (local_pf_num == 0 && local_vf_num == 934 && local_vf_active == 1) port_count[934]++; 
              else if (local_pf_num == 0 && local_vf_num == 935 && local_vf_active == 1) port_count[935]++; 
              else if (local_pf_num == 0 && local_vf_num == 936 && local_vf_active == 1) port_count[936]++; 
              else if (local_pf_num == 0 && local_vf_num == 937 && local_vf_active == 1) port_count[937]++; 
              else if (local_pf_num == 0 && local_vf_num == 938 && local_vf_active == 1) port_count[938]++; 
              else if (local_pf_num == 0 && local_vf_num == 939 && local_vf_active == 1) port_count[939]++; 
              else if (local_pf_num == 0 && local_vf_num == 940 && local_vf_active == 1) port_count[940]++; 
              else if (local_pf_num == 0 && local_vf_num == 941 && local_vf_active == 1) port_count[941]++; 
              else if (local_pf_num == 0 && local_vf_num == 942 && local_vf_active == 1) port_count[942]++; 
              else if (local_pf_num == 0 && local_vf_num == 943 && local_vf_active == 1) port_count[943]++; 
              else if (local_pf_num == 0 && local_vf_num == 944 && local_vf_active == 1) port_count[944]++; 
              else if (local_pf_num == 0 && local_vf_num == 945 && local_vf_active == 1) port_count[945]++; 
              else if (local_pf_num == 0 && local_vf_num == 946 && local_vf_active == 1) port_count[946]++; 
              else if (local_pf_num == 0 && local_vf_num == 947 && local_vf_active == 1) port_count[947]++; 
              else if (local_pf_num == 0 && local_vf_num == 948 && local_vf_active == 1) port_count[948]++; 
              else if (local_pf_num == 0 && local_vf_num == 949 && local_vf_active == 1) port_count[949]++; 
              else if (local_pf_num == 0 && local_vf_num == 950 && local_vf_active == 1) port_count[950]++; 
              else if (local_pf_num == 0 && local_vf_num == 951 && local_vf_active == 1) port_count[951]++; 
              else if (local_pf_num == 0 && local_vf_num == 952 && local_vf_active == 1) port_count[952]++; 
              else if (local_pf_num == 0 && local_vf_num == 953 && local_vf_active == 1) port_count[953]++; 
              else if (local_pf_num == 0 && local_vf_num == 954 && local_vf_active == 1) port_count[954]++; 
              else if (local_pf_num == 0 && local_vf_num == 955 && local_vf_active == 1) port_count[955]++; 
              else if (local_pf_num == 0 && local_vf_num == 956 && local_vf_active == 1) port_count[956]++; 
              else if (local_pf_num == 0 && local_vf_num == 957 && local_vf_active == 1) port_count[957]++; 
              else if (local_pf_num == 0 && local_vf_num == 958 && local_vf_active == 1) port_count[958]++; 
              else if (local_pf_num == 0 && local_vf_num == 959 && local_vf_active == 1) port_count[959]++; 
              else if (local_pf_num == 0 && local_vf_num == 960 && local_vf_active == 1) port_count[960]++; 
              else if (local_pf_num == 0 && local_vf_num == 961 && local_vf_active == 1) port_count[961]++; 
              else if (local_pf_num == 0 && local_vf_num == 962 && local_vf_active == 1) port_count[962]++; 
              else if (local_pf_num == 0 && local_vf_num == 963 && local_vf_active == 1) port_count[963]++; 
              else if (local_pf_num == 0 && local_vf_num == 964 && local_vf_active == 1) port_count[964]++; 
              else if (local_pf_num == 0 && local_vf_num == 965 && local_vf_active == 1) port_count[965]++; 
              else if (local_pf_num == 0 && local_vf_num == 966 && local_vf_active == 1) port_count[966]++; 
              else if (local_pf_num == 0 && local_vf_num == 967 && local_vf_active == 1) port_count[967]++; 
              else if (local_pf_num == 0 && local_vf_num == 968 && local_vf_active == 1) port_count[968]++; 
              else if (local_pf_num == 0 && local_vf_num == 969 && local_vf_active == 1) port_count[969]++; 
              else if (local_pf_num == 0 && local_vf_num == 970 && local_vf_active == 1) port_count[970]++; 
              else if (local_pf_num == 0 && local_vf_num == 971 && local_vf_active == 1) port_count[971]++; 
              else if (local_pf_num == 0 && local_vf_num == 972 && local_vf_active == 1) port_count[972]++; 
              else if (local_pf_num == 0 && local_vf_num == 973 && local_vf_active == 1) port_count[973]++; 
              else if (local_pf_num == 0 && local_vf_num == 974 && local_vf_active == 1) port_count[974]++; 
              else if (local_pf_num == 0 && local_vf_num == 975 && local_vf_active == 1) port_count[975]++; 
              else if (local_pf_num == 0 && local_vf_num == 976 && local_vf_active == 1) port_count[976]++; 
              else if (local_pf_num == 0 && local_vf_num == 977 && local_vf_active == 1) port_count[977]++; 
              else if (local_pf_num == 0 && local_vf_num == 978 && local_vf_active == 1) port_count[978]++; 
              else if (local_pf_num == 0 && local_vf_num == 979 && local_vf_active == 1) port_count[979]++; 
              else if (local_pf_num == 0 && local_vf_num == 980 && local_vf_active == 1) port_count[980]++; 
              else if (local_pf_num == 0 && local_vf_num == 981 && local_vf_active == 1) port_count[981]++; 
              else if (local_pf_num == 0 && local_vf_num == 982 && local_vf_active == 1) port_count[982]++; 
              else if (local_pf_num == 0 && local_vf_num == 983 && local_vf_active == 1) port_count[983]++; 
              else if (local_pf_num == 0 && local_vf_num == 984 && local_vf_active == 1) port_count[984]++; 
              else if (local_pf_num == 0 && local_vf_num == 985 && local_vf_active == 1) port_count[985]++; 
              else if (local_pf_num == 0 && local_vf_num == 986 && local_vf_active == 1) port_count[986]++; 
              else if (local_pf_num == 0 && local_vf_num == 987 && local_vf_active == 1) port_count[987]++; 
              else if (local_pf_num == 0 && local_vf_num == 988 && local_vf_active == 1) port_count[988]++; 
              else if (local_pf_num == 0 && local_vf_num == 989 && local_vf_active == 1) port_count[989]++; 
              else if (local_pf_num == 0 && local_vf_num == 990 && local_vf_active == 1) port_count[990]++; 
              else if (local_pf_num == 0 && local_vf_num == 991 && local_vf_active == 1) port_count[991]++; 
              else if (local_pf_num == 0 && local_vf_num == 992 && local_vf_active == 1) port_count[992]++; 
              else if (local_pf_num == 0 && local_vf_num == 993 && local_vf_active == 1) port_count[993]++; 
              else if (local_pf_num == 0 && local_vf_num == 994 && local_vf_active == 1) port_count[994]++; 
              else if (local_pf_num == 0 && local_vf_num == 995 && local_vf_active == 1) port_count[995]++; 
              else if (local_pf_num == 0 && local_vf_num == 996 && local_vf_active == 1) port_count[996]++; 
              else if (local_pf_num == 0 && local_vf_num == 997 && local_vf_active == 1) port_count[997]++; 
              else if (local_pf_num == 0 && local_vf_num == 998 && local_vf_active == 1) port_count[998]++; 
              else if (local_pf_num == 0 && local_vf_num == 999 && local_vf_active == 1) port_count[999]++; 
              else if (local_pf_num == 0 && local_vf_num == 1000 && local_vf_active == 1) port_count[1000]++; 
              else if (local_pf_num == 0 && local_vf_num == 1001 && local_vf_active == 1) port_count[1001]++; 
              else if (local_pf_num == 0 && local_vf_num == 1002 && local_vf_active == 1) port_count[1002]++; 
              else if (local_pf_num == 0 && local_vf_num == 1003 && local_vf_active == 1) port_count[1003]++; 
              else if (local_pf_num == 0 && local_vf_num == 1004 && local_vf_active == 1) port_count[1004]++; 
              else if (local_pf_num == 0 && local_vf_num == 1005 && local_vf_active == 1) port_count[1005]++; 
              else if (local_pf_num == 0 && local_vf_num == 1006 && local_vf_active == 1) port_count[1006]++; 
              else if (local_pf_num == 0 && local_vf_num == 1007 && local_vf_active == 1) port_count[1007]++; 
              else if (local_pf_num == 0 && local_vf_num == 1008 && local_vf_active == 1) port_count[1008]++; 
              else if (local_pf_num == 0 && local_vf_num == 1009 && local_vf_active == 1) port_count[1009]++; 
              else if (local_pf_num == 0 && local_vf_num == 1010 && local_vf_active == 1) port_count[1010]++; 
              else if (local_pf_num == 0 && local_vf_num == 1011 && local_vf_active == 1) port_count[1011]++; 
              else if (local_pf_num == 0 && local_vf_num == 1012 && local_vf_active == 1) port_count[1012]++; 
              else if (local_pf_num == 0 && local_vf_num == 1013 && local_vf_active == 1) port_count[1013]++; 
              else if (local_pf_num == 0 && local_vf_num == 1014 && local_vf_active == 1) port_count[1014]++; 
              else if (local_pf_num == 0 && local_vf_num == 1015 && local_vf_active == 1) port_count[1015]++; 
              else if (local_pf_num == 0 && local_vf_num == 1016 && local_vf_active == 1) port_count[1016]++; 
              else if (local_pf_num == 0 && local_vf_num == 1017 && local_vf_active == 1) port_count[1017]++; 
              else if (local_pf_num == 0 && local_vf_num == 1018 && local_vf_active == 1) port_count[1018]++; 
              else if (local_pf_num == 0 && local_vf_num == 1019 && local_vf_active == 1) port_count[1019]++; 
              else if (local_pf_num == 0 && local_vf_num == 1020 && local_vf_active == 1) port_count[1020]++; 
              else if (local_pf_num == 0 && local_vf_num == 1021 && local_vf_active == 1) port_count[1021]++; 
              else if (local_pf_num == 0 && local_vf_num == 1022 && local_vf_active == 1) port_count[1022]++; 
              else if (local_pf_num == 0 && local_vf_num == 1023 && local_vf_active == 1) port_count[1023]++; 
              else if (local_pf_num == 0 && local_vf_num == 1024 && local_vf_active == 1) port_count[1024]++; 
              else if (local_pf_num == 0 && local_vf_num == 1025 && local_vf_active == 1) port_count[1025]++; 
              else if (local_pf_num == 0 && local_vf_num == 1026 && local_vf_active == 1) port_count[1026]++; 
              else if (local_pf_num == 0 && local_vf_num == 1027 && local_vf_active == 1) port_count[1027]++; 
              else if (local_pf_num == 0 && local_vf_num == 1028 && local_vf_active == 1) port_count[1028]++; 
              else if (local_pf_num == 0 && local_vf_num == 1029 && local_vf_active == 1) port_count[1029]++; 
              else if (local_pf_num == 0 && local_vf_num == 1030 && local_vf_active == 1) port_count[1030]++; 
              else if (local_pf_num == 0 && local_vf_num == 1031 && local_vf_active == 1) port_count[1031]++; 
              else if (local_pf_num == 0 && local_vf_num == 1032 && local_vf_active == 1) port_count[1032]++; 
              else if (local_pf_num == 0 && local_vf_num == 1033 && local_vf_active == 1) port_count[1033]++; 
              else if (local_pf_num == 0 && local_vf_num == 1034 && local_vf_active == 1) port_count[1034]++; 
              else if (local_pf_num == 0 && local_vf_num == 1035 && local_vf_active == 1) port_count[1035]++; 
              else if (local_pf_num == 0 && local_vf_num == 1036 && local_vf_active == 1) port_count[1036]++; 
              else if (local_pf_num == 0 && local_vf_num == 1037 && local_vf_active == 1) port_count[1037]++; 
              else if (local_pf_num == 0 && local_vf_num == 1038 && local_vf_active == 1) port_count[1038]++; 
              else if (local_pf_num == 0 && local_vf_num == 1039 && local_vf_active == 1) port_count[1039]++; 
              else if (local_pf_num == 0 && local_vf_num == 1040 && local_vf_active == 1) port_count[1040]++; 
              else if (local_pf_num == 0 && local_vf_num == 1041 && local_vf_active == 1) port_count[1041]++; 
              else if (local_pf_num == 0 && local_vf_num == 1042 && local_vf_active == 1) port_count[1042]++; 
              else if (local_pf_num == 0 && local_vf_num == 1043 && local_vf_active == 1) port_count[1043]++; 
              else if (local_pf_num == 0 && local_vf_num == 1044 && local_vf_active == 1) port_count[1044]++; 
              else if (local_pf_num == 0 && local_vf_num == 1045 && local_vf_active == 1) port_count[1045]++; 
              else if (local_pf_num == 0 && local_vf_num == 1046 && local_vf_active == 1) port_count[1046]++; 
              else if (local_pf_num == 0 && local_vf_num == 1047 && local_vf_active == 1) port_count[1047]++; 
              else if (local_pf_num == 0 && local_vf_num == 1048 && local_vf_active == 1) port_count[1048]++; 
              else if (local_pf_num == 0 && local_vf_num == 1049 && local_vf_active == 1) port_count[1049]++; 
              else if (local_pf_num == 0 && local_vf_num == 1050 && local_vf_active == 1) port_count[1050]++; 
              else if (local_pf_num == 0 && local_vf_num == 1051 && local_vf_active == 1) port_count[1051]++; 
              else if (local_pf_num == 0 && local_vf_num == 1052 && local_vf_active == 1) port_count[1052]++; 
              else if (local_pf_num == 0 && local_vf_num == 1053 && local_vf_active == 1) port_count[1053]++; 
              else if (local_pf_num == 0 && local_vf_num == 1054 && local_vf_active == 1) port_count[1054]++; 
              else if (local_pf_num == 0 && local_vf_num == 1055 && local_vf_active == 1) port_count[1055]++; 
              else if (local_pf_num == 0 && local_vf_num == 1056 && local_vf_active == 1) port_count[1056]++; 
              else if (local_pf_num == 0 && local_vf_num == 1057 && local_vf_active == 1) port_count[1057]++; 
              else if (local_pf_num == 0 && local_vf_num == 1058 && local_vf_active == 1) port_count[1058]++; 
              else if (local_pf_num == 0 && local_vf_num == 1059 && local_vf_active == 1) port_count[1059]++; 
              else if (local_pf_num == 0 && local_vf_num == 1060 && local_vf_active == 1) port_count[1060]++; 
              else if (local_pf_num == 0 && local_vf_num == 1061 && local_vf_active == 1) port_count[1061]++; 
              else if (local_pf_num == 0 && local_vf_num == 1062 && local_vf_active == 1) port_count[1062]++; 
              else if (local_pf_num == 0 && local_vf_num == 1063 && local_vf_active == 1) port_count[1063]++; 
              else if (local_pf_num == 0 && local_vf_num == 1064 && local_vf_active == 1) port_count[1064]++; 
              else if (local_pf_num == 0 && local_vf_num == 1065 && local_vf_active == 1) port_count[1065]++; 
              else if (local_pf_num == 0 && local_vf_num == 1066 && local_vf_active == 1) port_count[1066]++; 
              else if (local_pf_num == 0 && local_vf_num == 1067 && local_vf_active == 1) port_count[1067]++; 
              else if (local_pf_num == 0 && local_vf_num == 1068 && local_vf_active == 1) port_count[1068]++; 
              else if (local_pf_num == 0 && local_vf_num == 1069 && local_vf_active == 1) port_count[1069]++; 
              else if (local_pf_num == 0 && local_vf_num == 1070 && local_vf_active == 1) port_count[1070]++; 
              else if (local_pf_num == 0 && local_vf_num == 1071 && local_vf_active == 1) port_count[1071]++; 
              else if (local_pf_num == 0 && local_vf_num == 1072 && local_vf_active == 1) port_count[1072]++; 
              else if (local_pf_num == 0 && local_vf_num == 1073 && local_vf_active == 1) port_count[1073]++; 
              else if (local_pf_num == 0 && local_vf_num == 1074 && local_vf_active == 1) port_count[1074]++; 
              else if (local_pf_num == 0 && local_vf_num == 1075 && local_vf_active == 1) port_count[1075]++; 
              else if (local_pf_num == 0 && local_vf_num == 1076 && local_vf_active == 1) port_count[1076]++; 
              else if (local_pf_num == 0 && local_vf_num == 1077 && local_vf_active == 1) port_count[1077]++; 
              else if (local_pf_num == 0 && local_vf_num == 1078 && local_vf_active == 1) port_count[1078]++; 
              else if (local_pf_num == 0 && local_vf_num == 1079 && local_vf_active == 1) port_count[1079]++; 
              else if (local_pf_num == 0 && local_vf_num == 1080 && local_vf_active == 1) port_count[1080]++; 
              else if (local_pf_num == 0 && local_vf_num == 1081 && local_vf_active == 1) port_count[1081]++; 
              else if (local_pf_num == 0 && local_vf_num == 1082 && local_vf_active == 1) port_count[1082]++; 
              else if (local_pf_num == 0 && local_vf_num == 1083 && local_vf_active == 1) port_count[1083]++; 
              else if (local_pf_num == 0 && local_vf_num == 1084 && local_vf_active == 1) port_count[1084]++; 
              else if (local_pf_num == 0 && local_vf_num == 1085 && local_vf_active == 1) port_count[1085]++; 
              else if (local_pf_num == 0 && local_vf_num == 1086 && local_vf_active == 1) port_count[1086]++; 
              else if (local_pf_num == 0 && local_vf_num == 1087 && local_vf_active == 1) port_count[1087]++; 
              else if (local_pf_num == 0 && local_vf_num == 1088 && local_vf_active == 1) port_count[1088]++; 
              else if (local_pf_num == 0 && local_vf_num == 1089 && local_vf_active == 1) port_count[1089]++; 
              else if (local_pf_num == 0 && local_vf_num == 1090 && local_vf_active == 1) port_count[1090]++; 
              else if (local_pf_num == 0 && local_vf_num == 1091 && local_vf_active == 1) port_count[1091]++; 
              else if (local_pf_num == 0 && local_vf_num == 1092 && local_vf_active == 1) port_count[1092]++; 
              else if (local_pf_num == 0 && local_vf_num == 1093 && local_vf_active == 1) port_count[1093]++; 
              else if (local_pf_num == 0 && local_vf_num == 1094 && local_vf_active == 1) port_count[1094]++; 
              else if (local_pf_num == 0 && local_vf_num == 1095 && local_vf_active == 1) port_count[1095]++; 
              else if (local_pf_num == 0 && local_vf_num == 1096 && local_vf_active == 1) port_count[1096]++; 
              else if (local_pf_num == 0 && local_vf_num == 1097 && local_vf_active == 1) port_count[1097]++; 
              else if (local_pf_num == 0 && local_vf_num == 1098 && local_vf_active == 1) port_count[1098]++; 
              else if (local_pf_num == 0 && local_vf_num == 1099 && local_vf_active == 1) port_count[1099]++; 
              else if (local_pf_num == 0 && local_vf_num == 1100 && local_vf_active == 1) port_count[1100]++; 
              else if (local_pf_num == 0 && local_vf_num == 1101 && local_vf_active == 1) port_count[1101]++; 
              else if (local_pf_num == 0 && local_vf_num == 1102 && local_vf_active == 1) port_count[1102]++; 
              else if (local_pf_num == 0 && local_vf_num == 1103 && local_vf_active == 1) port_count[1103]++; 
              else if (local_pf_num == 0 && local_vf_num == 1104 && local_vf_active == 1) port_count[1104]++; 
              else if (local_pf_num == 0 && local_vf_num == 1105 && local_vf_active == 1) port_count[1105]++; 
              else if (local_pf_num == 0 && local_vf_num == 1106 && local_vf_active == 1) port_count[1106]++; 
              else if (local_pf_num == 0 && local_vf_num == 1107 && local_vf_active == 1) port_count[1107]++; 
              else if (local_pf_num == 0 && local_vf_num == 1108 && local_vf_active == 1) port_count[1108]++; 
              else if (local_pf_num == 0 && local_vf_num == 1109 && local_vf_active == 1) port_count[1109]++; 
              else if (local_pf_num == 0 && local_vf_num == 1110 && local_vf_active == 1) port_count[1110]++; 
              else if (local_pf_num == 0 && local_vf_num == 1111 && local_vf_active == 1) port_count[1111]++; 
              else if (local_pf_num == 0 && local_vf_num == 1112 && local_vf_active == 1) port_count[1112]++; 
              else if (local_pf_num == 0 && local_vf_num == 1113 && local_vf_active == 1) port_count[1113]++; 
              else if (local_pf_num == 0 && local_vf_num == 1114 && local_vf_active == 1) port_count[1114]++; 
              else if (local_pf_num == 0 && local_vf_num == 1115 && local_vf_active == 1) port_count[1115]++; 
              else if (local_pf_num == 0 && local_vf_num == 1116 && local_vf_active == 1) port_count[1116]++; 
              else if (local_pf_num == 0 && local_vf_num == 1117 && local_vf_active == 1) port_count[1117]++; 
              else if (local_pf_num == 0 && local_vf_num == 1118 && local_vf_active == 1) port_count[1118]++; 
              else if (local_pf_num == 0 && local_vf_num == 1119 && local_vf_active == 1) port_count[1119]++; 
              else if (local_pf_num == 0 && local_vf_num == 1120 && local_vf_active == 1) port_count[1120]++; 
              else if (local_pf_num == 0 && local_vf_num == 1121 && local_vf_active == 1) port_count[1121]++; 
              else if (local_pf_num == 0 && local_vf_num == 1122 && local_vf_active == 1) port_count[1122]++; 
              else if (local_pf_num == 0 && local_vf_num == 1123 && local_vf_active == 1) port_count[1123]++; 
              else if (local_pf_num == 0 && local_vf_num == 1124 && local_vf_active == 1) port_count[1124]++; 
              else if (local_pf_num == 0 && local_vf_num == 1125 && local_vf_active == 1) port_count[1125]++; 
              else if (local_pf_num == 0 && local_vf_num == 1126 && local_vf_active == 1) port_count[1126]++; 
              else if (local_pf_num == 0 && local_vf_num == 1127 && local_vf_active == 1) port_count[1127]++; 
              else if (local_pf_num == 0 && local_vf_num == 1128 && local_vf_active == 1) port_count[1128]++; 
              else if (local_pf_num == 0 && local_vf_num == 1129 && local_vf_active == 1) port_count[1129]++; 
              else if (local_pf_num == 0 && local_vf_num == 1130 && local_vf_active == 1) port_count[1130]++; 
              else if (local_pf_num == 0 && local_vf_num == 1131 && local_vf_active == 1) port_count[1131]++; 
              else if (local_pf_num == 0 && local_vf_num == 1132 && local_vf_active == 1) port_count[1132]++; 
              else if (local_pf_num == 0 && local_vf_num == 1133 && local_vf_active == 1) port_count[1133]++; 
              else if (local_pf_num == 0 && local_vf_num == 1134 && local_vf_active == 1) port_count[1134]++; 
              else if (local_pf_num == 0 && local_vf_num == 1135 && local_vf_active == 1) port_count[1135]++; 
              else if (local_pf_num == 0 && local_vf_num == 1136 && local_vf_active == 1) port_count[1136]++; 
              else if (local_pf_num == 0 && local_vf_num == 1137 && local_vf_active == 1) port_count[1137]++; 
              else if (local_pf_num == 0 && local_vf_num == 1138 && local_vf_active == 1) port_count[1138]++; 
              else if (local_pf_num == 0 && local_vf_num == 1139 && local_vf_active == 1) port_count[1139]++; 
              else if (local_pf_num == 0 && local_vf_num == 1140 && local_vf_active == 1) port_count[1140]++; 
              else if (local_pf_num == 0 && local_vf_num == 1141 && local_vf_active == 1) port_count[1141]++; 
              else if (local_pf_num == 0 && local_vf_num == 1142 && local_vf_active == 1) port_count[1142]++; 
              else if (local_pf_num == 0 && local_vf_num == 1143 && local_vf_active == 1) port_count[1143]++; 
              else if (local_pf_num == 0 && local_vf_num == 1144 && local_vf_active == 1) port_count[1144]++; 
              else if (local_pf_num == 0 && local_vf_num == 1145 && local_vf_active == 1) port_count[1145]++; 
              else if (local_pf_num == 0 && local_vf_num == 1146 && local_vf_active == 1) port_count[1146]++; 
              else if (local_pf_num == 0 && local_vf_num == 1147 && local_vf_active == 1) port_count[1147]++; 
              else if (local_pf_num == 0 && local_vf_num == 1148 && local_vf_active == 1) port_count[1148]++; 
              else if (local_pf_num == 0 && local_vf_num == 1149 && local_vf_active == 1) port_count[1149]++; 
              else if (local_pf_num == 0 && local_vf_num == 1150 && local_vf_active == 1) port_count[1150]++; 
              else if (local_pf_num == 0 && local_vf_num == 1151 && local_vf_active == 1) port_count[1151]++; 
              else if (local_pf_num == 0 && local_vf_num == 1152 && local_vf_active == 1) port_count[1152]++; 
              else if (local_pf_num == 0 && local_vf_num == 1153 && local_vf_active == 1) port_count[1153]++; 
              else if (local_pf_num == 0 && local_vf_num == 1154 && local_vf_active == 1) port_count[1154]++; 
              else if (local_pf_num == 0 && local_vf_num == 1155 && local_vf_active == 1) port_count[1155]++; 
              else if (local_pf_num == 0 && local_vf_num == 1156 && local_vf_active == 1) port_count[1156]++; 
              else if (local_pf_num == 0 && local_vf_num == 1157 && local_vf_active == 1) port_count[1157]++; 
              else if (local_pf_num == 0 && local_vf_num == 1158 && local_vf_active == 1) port_count[1158]++; 
              else if (local_pf_num == 0 && local_vf_num == 1159 && local_vf_active == 1) port_count[1159]++; 
              else if (local_pf_num == 0 && local_vf_num == 1160 && local_vf_active == 1) port_count[1160]++; 
              else if (local_pf_num == 0 && local_vf_num == 1161 && local_vf_active == 1) port_count[1161]++; 
              else if (local_pf_num == 0 && local_vf_num == 1162 && local_vf_active == 1) port_count[1162]++; 
              else if (local_pf_num == 0 && local_vf_num == 1163 && local_vf_active == 1) port_count[1163]++; 
              else if (local_pf_num == 0 && local_vf_num == 1164 && local_vf_active == 1) port_count[1164]++; 
              else if (local_pf_num == 0 && local_vf_num == 1165 && local_vf_active == 1) port_count[1165]++; 
              else if (local_pf_num == 0 && local_vf_num == 1166 && local_vf_active == 1) port_count[1166]++; 
              else if (local_pf_num == 0 && local_vf_num == 1167 && local_vf_active == 1) port_count[1167]++; 
              else if (local_pf_num == 0 && local_vf_num == 1168 && local_vf_active == 1) port_count[1168]++; 
              else if (local_pf_num == 0 && local_vf_num == 1169 && local_vf_active == 1) port_count[1169]++; 
              else if (local_pf_num == 0 && local_vf_num == 1170 && local_vf_active == 1) port_count[1170]++; 
              else if (local_pf_num == 0 && local_vf_num == 1171 && local_vf_active == 1) port_count[1171]++; 
              else if (local_pf_num == 0 && local_vf_num == 1172 && local_vf_active == 1) port_count[1172]++; 
              else if (local_pf_num == 0 && local_vf_num == 1173 && local_vf_active == 1) port_count[1173]++; 
              else if (local_pf_num == 0 && local_vf_num == 1174 && local_vf_active == 1) port_count[1174]++; 
              else if (local_pf_num == 0 && local_vf_num == 1175 && local_vf_active == 1) port_count[1175]++; 
              else if (local_pf_num == 0 && local_vf_num == 1176 && local_vf_active == 1) port_count[1176]++; 
              else if (local_pf_num == 0 && local_vf_num == 1177 && local_vf_active == 1) port_count[1177]++; 
              else if (local_pf_num == 0 && local_vf_num == 1178 && local_vf_active == 1) port_count[1178]++; 
              else if (local_pf_num == 0 && local_vf_num == 1179 && local_vf_active == 1) port_count[1179]++; 
              else if (local_pf_num == 0 && local_vf_num == 1180 && local_vf_active == 1) port_count[1180]++; 
              else if (local_pf_num == 0 && local_vf_num == 1181 && local_vf_active == 1) port_count[1181]++; 
              else if (local_pf_num == 0 && local_vf_num == 1182 && local_vf_active == 1) port_count[1182]++; 
              else if (local_pf_num == 0 && local_vf_num == 1183 && local_vf_active == 1) port_count[1183]++; 
              else if (local_pf_num == 0 && local_vf_num == 1184 && local_vf_active == 1) port_count[1184]++; 
              else if (local_pf_num == 0 && local_vf_num == 1185 && local_vf_active == 1) port_count[1185]++; 
              else if (local_pf_num == 0 && local_vf_num == 1186 && local_vf_active == 1) port_count[1186]++; 
              else if (local_pf_num == 0 && local_vf_num == 1187 && local_vf_active == 1) port_count[1187]++; 
              else if (local_pf_num == 0 && local_vf_num == 1188 && local_vf_active == 1) port_count[1188]++; 
              else if (local_pf_num == 0 && local_vf_num == 1189 && local_vf_active == 1) port_count[1189]++; 
              else if (local_pf_num == 0 && local_vf_num == 1190 && local_vf_active == 1) port_count[1190]++; 
              else if (local_pf_num == 0 && local_vf_num == 1191 && local_vf_active == 1) port_count[1191]++; 
              else if (local_pf_num == 0 && local_vf_num == 1192 && local_vf_active == 1) port_count[1192]++; 
              else if (local_pf_num == 0 && local_vf_num == 1193 && local_vf_active == 1) port_count[1193]++; 
              else if (local_pf_num == 0 && local_vf_num == 1194 && local_vf_active == 1) port_count[1194]++; 
              else if (local_pf_num == 0 && local_vf_num == 1195 && local_vf_active == 1) port_count[1195]++; 
              else if (local_pf_num == 0 && local_vf_num == 1196 && local_vf_active == 1) port_count[1196]++; 
              else if (local_pf_num == 0 && local_vf_num == 1197 && local_vf_active == 1) port_count[1197]++; 
              else if (local_pf_num == 0 && local_vf_num == 1198 && local_vf_active == 1) port_count[1198]++; 
              else if (local_pf_num == 0 && local_vf_num == 1199 && local_vf_active == 1) port_count[1199]++; 
              else if (local_pf_num == 0 && local_vf_num == 1200 && local_vf_active == 1) port_count[1200]++; 
              else if (local_pf_num == 0 && local_vf_num == 1201 && local_vf_active == 1) port_count[1201]++; 
              else if (local_pf_num == 0 && local_vf_num == 1202 && local_vf_active == 1) port_count[1202]++; 
              else if (local_pf_num == 0 && local_vf_num == 1203 && local_vf_active == 1) port_count[1203]++; 
              else if (local_pf_num == 0 && local_vf_num == 1204 && local_vf_active == 1) port_count[1204]++; 
              else if (local_pf_num == 0 && local_vf_num == 1205 && local_vf_active == 1) port_count[1205]++; 
              else if (local_pf_num == 0 && local_vf_num == 1206 && local_vf_active == 1) port_count[1206]++; 
              else if (local_pf_num == 0 && local_vf_num == 1207 && local_vf_active == 1) port_count[1207]++; 
              else if (local_pf_num == 0 && local_vf_num == 1208 && local_vf_active == 1) port_count[1208]++; 
              else if (local_pf_num == 0 && local_vf_num == 1209 && local_vf_active == 1) port_count[1209]++; 
              else if (local_pf_num == 0 && local_vf_num == 1210 && local_vf_active == 1) port_count[1210]++; 
              else if (local_pf_num == 0 && local_vf_num == 1211 && local_vf_active == 1) port_count[1211]++; 
              else if (local_pf_num == 0 && local_vf_num == 1212 && local_vf_active == 1) port_count[1212]++; 
              else if (local_pf_num == 0 && local_vf_num == 1213 && local_vf_active == 1) port_count[1213]++; 
              else if (local_pf_num == 0 && local_vf_num == 1214 && local_vf_active == 1) port_count[1214]++; 
              else if (local_pf_num == 0 && local_vf_num == 1215 && local_vf_active == 1) port_count[1215]++; 
              else if (local_pf_num == 0 && local_vf_num == 1216 && local_vf_active == 1) port_count[1216]++; 
              else if (local_pf_num == 0 && local_vf_num == 1217 && local_vf_active == 1) port_count[1217]++; 
              else if (local_pf_num == 0 && local_vf_num == 1218 && local_vf_active == 1) port_count[1218]++; 
              else if (local_pf_num == 0 && local_vf_num == 1219 && local_vf_active == 1) port_count[1219]++; 
              else if (local_pf_num == 0 && local_vf_num == 1220 && local_vf_active == 1) port_count[1220]++; 
              else if (local_pf_num == 0 && local_vf_num == 1221 && local_vf_active == 1) port_count[1221]++; 
              else if (local_pf_num == 0 && local_vf_num == 1222 && local_vf_active == 1) port_count[1222]++; 
              else if (local_pf_num == 0 && local_vf_num == 1223 && local_vf_active == 1) port_count[1223]++; 
              else if (local_pf_num == 0 && local_vf_num == 1224 && local_vf_active == 1) port_count[1224]++; 
              else if (local_pf_num == 0 && local_vf_num == 1225 && local_vf_active == 1) port_count[1225]++; 
              else if (local_pf_num == 0 && local_vf_num == 1226 && local_vf_active == 1) port_count[1226]++; 
              else if (local_pf_num == 0 && local_vf_num == 1227 && local_vf_active == 1) port_count[1227]++; 
              else if (local_pf_num == 0 && local_vf_num == 1228 && local_vf_active == 1) port_count[1228]++; 
              else if (local_pf_num == 0 && local_vf_num == 1229 && local_vf_active == 1) port_count[1229]++; 
              else if (local_pf_num == 0 && local_vf_num == 1230 && local_vf_active == 1) port_count[1230]++; 
              else if (local_pf_num == 0 && local_vf_num == 1231 && local_vf_active == 1) port_count[1231]++; 
              else if (local_pf_num == 0 && local_vf_num == 1232 && local_vf_active == 1) port_count[1232]++; 
              else if (local_pf_num == 0 && local_vf_num == 1233 && local_vf_active == 1) port_count[1233]++; 
              else if (local_pf_num == 0 && local_vf_num == 1234 && local_vf_active == 1) port_count[1234]++; 
              else if (local_pf_num == 0 && local_vf_num == 1235 && local_vf_active == 1) port_count[1235]++; 
              else if (local_pf_num == 0 && local_vf_num == 1236 && local_vf_active == 1) port_count[1236]++; 
              else if (local_pf_num == 0 && local_vf_num == 1237 && local_vf_active == 1) port_count[1237]++; 
              else if (local_pf_num == 0 && local_vf_num == 1238 && local_vf_active == 1) port_count[1238]++; 
              else if (local_pf_num == 0 && local_vf_num == 1239 && local_vf_active == 1) port_count[1239]++; 
              else if (local_pf_num == 0 && local_vf_num == 1240 && local_vf_active == 1) port_count[1240]++; 
              else if (local_pf_num == 0 && local_vf_num == 1241 && local_vf_active == 1) port_count[1241]++; 
              else if (local_pf_num == 0 && local_vf_num == 1242 && local_vf_active == 1) port_count[1242]++; 
              else if (local_pf_num == 0 && local_vf_num == 1243 && local_vf_active == 1) port_count[1243]++; 
              else if (local_pf_num == 0 && local_vf_num == 1244 && local_vf_active == 1) port_count[1244]++; 
              else if (local_pf_num == 0 && local_vf_num == 1245 && local_vf_active == 1) port_count[1245]++; 
              else if (local_pf_num == 0 && local_vf_num == 1246 && local_vf_active == 1) port_count[1246]++; 
              else if (local_pf_num == 0 && local_vf_num == 1247 && local_vf_active == 1) port_count[1247]++; 
              else if (local_pf_num == 0 && local_vf_num == 1248 && local_vf_active == 1) port_count[1248]++; 
              else if (local_pf_num == 0 && local_vf_num == 1249 && local_vf_active == 1) port_count[1249]++; 
              else if (local_pf_num == 0 && local_vf_num == 1250 && local_vf_active == 1) port_count[1250]++; 
              else if (local_pf_num == 0 && local_vf_num == 1251 && local_vf_active == 1) port_count[1251]++; 
              else if (local_pf_num == 0 && local_vf_num == 1252 && local_vf_active == 1) port_count[1252]++; 
              else if (local_pf_num == 0 && local_vf_num == 1253 && local_vf_active == 1) port_count[1253]++; 
              else if (local_pf_num == 0 && local_vf_num == 1254 && local_vf_active == 1) port_count[1254]++; 
              else if (local_pf_num == 0 && local_vf_num == 1255 && local_vf_active == 1) port_count[1255]++; 
              else if (local_pf_num == 0 && local_vf_num == 1256 && local_vf_active == 1) port_count[1256]++; 
              else if (local_pf_num == 0 && local_vf_num == 1257 && local_vf_active == 1) port_count[1257]++; 
              else if (local_pf_num == 0 && local_vf_num == 1258 && local_vf_active == 1) port_count[1258]++; 
              else if (local_pf_num == 0 && local_vf_num == 1259 && local_vf_active == 1) port_count[1259]++; 
              else if (local_pf_num == 0 && local_vf_num == 1260 && local_vf_active == 1) port_count[1260]++; 
              else if (local_pf_num == 0 && local_vf_num == 1261 && local_vf_active == 1) port_count[1261]++; 
              else if (local_pf_num == 0 && local_vf_num == 1262 && local_vf_active == 1) port_count[1262]++; 
              else if (local_pf_num == 0 && local_vf_num == 1263 && local_vf_active == 1) port_count[1263]++; 
              else if (local_pf_num == 0 && local_vf_num == 1264 && local_vf_active == 1) port_count[1264]++; 
              else if (local_pf_num == 0 && local_vf_num == 1265 && local_vf_active == 1) port_count[1265]++; 
              else if (local_pf_num == 0 && local_vf_num == 1266 && local_vf_active == 1) port_count[1266]++; 
              else if (local_pf_num == 0 && local_vf_num == 1267 && local_vf_active == 1) port_count[1267]++; 
              else if (local_pf_num == 0 && local_vf_num == 1268 && local_vf_active == 1) port_count[1268]++; 
              else if (local_pf_num == 0 && local_vf_num == 1269 && local_vf_active == 1) port_count[1269]++; 
              else if (local_pf_num == 0 && local_vf_num == 1270 && local_vf_active == 1) port_count[1270]++; 
              else if (local_pf_num == 0 && local_vf_num == 1271 && local_vf_active == 1) port_count[1271]++; 
              else if (local_pf_num == 0 && local_vf_num == 1272 && local_vf_active == 1) port_count[1272]++; 
              else if (local_pf_num == 0 && local_vf_num == 1273 && local_vf_active == 1) port_count[1273]++; 
              else if (local_pf_num == 0 && local_vf_num == 1274 && local_vf_active == 1) port_count[1274]++; 
              else if (local_pf_num == 0 && local_vf_num == 1275 && local_vf_active == 1) port_count[1275]++; 
              else if (local_pf_num == 0 && local_vf_num == 1276 && local_vf_active == 1) port_count[1276]++; 
              else if (local_pf_num == 0 && local_vf_num == 1277 && local_vf_active == 1) port_count[1277]++; 
              else if (local_pf_num == 0 && local_vf_num == 1278 && local_vf_active == 1) port_count[1278]++; 
              else if (local_pf_num == 0 && local_vf_num == 1279 && local_vf_active == 1) port_count[1279]++; 
              else if (local_pf_num == 0 && local_vf_num == 1280 && local_vf_active == 1) port_count[1280]++; 
              else if (local_pf_num == 0 && local_vf_num == 1281 && local_vf_active == 1) port_count[1281]++; 
              else if (local_pf_num == 0 && local_vf_num == 1282 && local_vf_active == 1) port_count[1282]++; 
              else if (local_pf_num == 0 && local_vf_num == 1283 && local_vf_active == 1) port_count[1283]++; 
              else if (local_pf_num == 0 && local_vf_num == 1284 && local_vf_active == 1) port_count[1284]++; 
              else if (local_pf_num == 0 && local_vf_num == 1285 && local_vf_active == 1) port_count[1285]++; 
              else if (local_pf_num == 0 && local_vf_num == 1286 && local_vf_active == 1) port_count[1286]++; 
              else if (local_pf_num == 0 && local_vf_num == 1287 && local_vf_active == 1) port_count[1287]++; 
              else if (local_pf_num == 0 && local_vf_num == 1288 && local_vf_active == 1) port_count[1288]++; 
              else if (local_pf_num == 0 && local_vf_num == 1289 && local_vf_active == 1) port_count[1289]++; 
              else if (local_pf_num == 0 && local_vf_num == 1290 && local_vf_active == 1) port_count[1290]++; 
              else if (local_pf_num == 0 && local_vf_num == 1291 && local_vf_active == 1) port_count[1291]++; 
              else if (local_pf_num == 0 && local_vf_num == 1292 && local_vf_active == 1) port_count[1292]++; 
              else if (local_pf_num == 0 && local_vf_num == 1293 && local_vf_active == 1) port_count[1293]++; 
              else if (local_pf_num == 0 && local_vf_num == 1294 && local_vf_active == 1) port_count[1294]++; 
              else if (local_pf_num == 0 && local_vf_num == 1295 && local_vf_active == 1) port_count[1295]++; 
              else if (local_pf_num == 0 && local_vf_num == 1296 && local_vf_active == 1) port_count[1296]++; 
              else if (local_pf_num == 0 && local_vf_num == 1297 && local_vf_active == 1) port_count[1297]++; 
              else if (local_pf_num == 0 && local_vf_num == 1298 && local_vf_active == 1) port_count[1298]++; 
              else if (local_pf_num == 0 && local_vf_num == 1299 && local_vf_active == 1) port_count[1299]++; 
              else if (local_pf_num == 0 && local_vf_num == 1300 && local_vf_active == 1) port_count[1300]++; 
              else if (local_pf_num == 0 && local_vf_num == 1301 && local_vf_active == 1) port_count[1301]++; 
              else if (local_pf_num == 0 && local_vf_num == 1302 && local_vf_active == 1) port_count[1302]++; 
              else if (local_pf_num == 0 && local_vf_num == 1303 && local_vf_active == 1) port_count[1303]++; 
              else if (local_pf_num == 0 && local_vf_num == 1304 && local_vf_active == 1) port_count[1304]++; 
              else if (local_pf_num == 0 && local_vf_num == 1305 && local_vf_active == 1) port_count[1305]++; 
              else if (local_pf_num == 0 && local_vf_num == 1306 && local_vf_active == 1) port_count[1306]++; 
              else if (local_pf_num == 0 && local_vf_num == 1307 && local_vf_active == 1) port_count[1307]++; 
              else if (local_pf_num == 0 && local_vf_num == 1308 && local_vf_active == 1) port_count[1308]++; 
              else if (local_pf_num == 0 && local_vf_num == 1309 && local_vf_active == 1) port_count[1309]++; 
              else if (local_pf_num == 0 && local_vf_num == 1310 && local_vf_active == 1) port_count[1310]++; 
              else if (local_pf_num == 0 && local_vf_num == 1311 && local_vf_active == 1) port_count[1311]++; 
              else if (local_pf_num == 0 && local_vf_num == 1312 && local_vf_active == 1) port_count[1312]++; 
              else if (local_pf_num == 0 && local_vf_num == 1313 && local_vf_active == 1) port_count[1313]++; 
              else if (local_pf_num == 0 && local_vf_num == 1314 && local_vf_active == 1) port_count[1314]++; 
              else if (local_pf_num == 0 && local_vf_num == 1315 && local_vf_active == 1) port_count[1315]++; 
              else if (local_pf_num == 0 && local_vf_num == 1316 && local_vf_active == 1) port_count[1316]++; 
              else if (local_pf_num == 0 && local_vf_num == 1317 && local_vf_active == 1) port_count[1317]++; 
              else if (local_pf_num == 0 && local_vf_num == 1318 && local_vf_active == 1) port_count[1318]++; 
              else if (local_pf_num == 0 && local_vf_num == 1319 && local_vf_active == 1) port_count[1319]++; 
              else if (local_pf_num == 0 && local_vf_num == 1320 && local_vf_active == 1) port_count[1320]++; 
              else if (local_pf_num == 0 && local_vf_num == 1321 && local_vf_active == 1) port_count[1321]++; 
              else if (local_pf_num == 0 && local_vf_num == 1322 && local_vf_active == 1) port_count[1322]++; 
              else if (local_pf_num == 0 && local_vf_num == 1323 && local_vf_active == 1) port_count[1323]++; 
              else if (local_pf_num == 0 && local_vf_num == 1324 && local_vf_active == 1) port_count[1324]++; 
              else if (local_pf_num == 0 && local_vf_num == 1325 && local_vf_active == 1) port_count[1325]++; 
              else if (local_pf_num == 0 && local_vf_num == 1326 && local_vf_active == 1) port_count[1326]++; 
              else if (local_pf_num == 0 && local_vf_num == 1327 && local_vf_active == 1) port_count[1327]++; 
              else if (local_pf_num == 0 && local_vf_num == 1328 && local_vf_active == 1) port_count[1328]++; 
              else if (local_pf_num == 0 && local_vf_num == 1329 && local_vf_active == 1) port_count[1329]++; 
              else if (local_pf_num == 0 && local_vf_num == 1330 && local_vf_active == 1) port_count[1330]++; 
              else if (local_pf_num == 0 && local_vf_num == 1331 && local_vf_active == 1) port_count[1331]++; 
              else if (local_pf_num == 0 && local_vf_num == 1332 && local_vf_active == 1) port_count[1332]++; 
              else if (local_pf_num == 0 && local_vf_num == 1333 && local_vf_active == 1) port_count[1333]++; 
              else if (local_pf_num == 0 && local_vf_num == 1334 && local_vf_active == 1) port_count[1334]++; 
              else if (local_pf_num == 0 && local_vf_num == 1335 && local_vf_active == 1) port_count[1335]++; 
              else if (local_pf_num == 0 && local_vf_num == 1336 && local_vf_active == 1) port_count[1336]++; 
              else if (local_pf_num == 0 && local_vf_num == 1337 && local_vf_active == 1) port_count[1337]++; 
              else if (local_pf_num == 0 && local_vf_num == 1338 && local_vf_active == 1) port_count[1338]++; 
              else if (local_pf_num == 0 && local_vf_num == 1339 && local_vf_active == 1) port_count[1339]++; 
              else if (local_pf_num == 0 && local_vf_num == 1340 && local_vf_active == 1) port_count[1340]++; 
              else if (local_pf_num == 0 && local_vf_num == 1341 && local_vf_active == 1) port_count[1341]++; 
              else if (local_pf_num == 0 && local_vf_num == 1342 && local_vf_active == 1) port_count[1342]++; 
              else if (local_pf_num == 0 && local_vf_num == 1343 && local_vf_active == 1) port_count[1343]++; 
              else if (local_pf_num == 0 && local_vf_num == 1344 && local_vf_active == 1) port_count[1344]++; 
              else if (local_pf_num == 0 && local_vf_num == 1345 && local_vf_active == 1) port_count[1345]++; 
              else if (local_pf_num == 0 && local_vf_num == 1346 && local_vf_active == 1) port_count[1346]++; 
              else if (local_pf_num == 0 && local_vf_num == 1347 && local_vf_active == 1) port_count[1347]++; 
              else if (local_pf_num == 0 && local_vf_num == 1348 && local_vf_active == 1) port_count[1348]++; 
              else if (local_pf_num == 0 && local_vf_num == 1349 && local_vf_active == 1) port_count[1349]++; 
              else if (local_pf_num == 0 && local_vf_num == 1350 && local_vf_active == 1) port_count[1350]++; 
              else if (local_pf_num == 0 && local_vf_num == 1351 && local_vf_active == 1) port_count[1351]++; 
              else if (local_pf_num == 0 && local_vf_num == 1352 && local_vf_active == 1) port_count[1352]++; 
              else if (local_pf_num == 0 && local_vf_num == 1353 && local_vf_active == 1) port_count[1353]++; 
              else if (local_pf_num == 0 && local_vf_num == 1354 && local_vf_active == 1) port_count[1354]++; 
              else if (local_pf_num == 0 && local_vf_num == 1355 && local_vf_active == 1) port_count[1355]++; 
              else if (local_pf_num == 0 && local_vf_num == 1356 && local_vf_active == 1) port_count[1356]++; 
              else if (local_pf_num == 0 && local_vf_num == 1357 && local_vf_active == 1) port_count[1357]++; 
              else if (local_pf_num == 0 && local_vf_num == 1358 && local_vf_active == 1) port_count[1358]++; 
              else if (local_pf_num == 0 && local_vf_num == 1359 && local_vf_active == 1) port_count[1359]++; 
              else if (local_pf_num == 0 && local_vf_num == 1360 && local_vf_active == 1) port_count[1360]++; 
              else if (local_pf_num == 0 && local_vf_num == 1361 && local_vf_active == 1) port_count[1361]++; 
              else if (local_pf_num == 0 && local_vf_num == 1362 && local_vf_active == 1) port_count[1362]++; 
              else if (local_pf_num == 0 && local_vf_num == 1363 && local_vf_active == 1) port_count[1363]++; 
              else if (local_pf_num == 0 && local_vf_num == 1364 && local_vf_active == 1) port_count[1364]++; 
              else if (local_pf_num == 0 && local_vf_num == 1365 && local_vf_active == 1) port_count[1365]++; 
              else if (local_pf_num == 0 && local_vf_num == 1366 && local_vf_active == 1) port_count[1366]++; 
              else if (local_pf_num == 0 && local_vf_num == 1367 && local_vf_active == 1) port_count[1367]++; 
              else if (local_pf_num == 0 && local_vf_num == 1368 && local_vf_active == 1) port_count[1368]++; 
              else if (local_pf_num == 0 && local_vf_num == 1369 && local_vf_active == 1) port_count[1369]++; 
              else if (local_pf_num == 0 && local_vf_num == 1370 && local_vf_active == 1) port_count[1370]++; 
              else if (local_pf_num == 0 && local_vf_num == 1371 && local_vf_active == 1) port_count[1371]++; 
              else if (local_pf_num == 0 && local_vf_num == 1372 && local_vf_active == 1) port_count[1372]++; 
              else if (local_pf_num == 0 && local_vf_num == 1373 && local_vf_active == 1) port_count[1373]++; 
              else if (local_pf_num == 0 && local_vf_num == 1374 && local_vf_active == 1) port_count[1374]++; 
              else if (local_pf_num == 0 && local_vf_num == 1375 && local_vf_active == 1) port_count[1375]++; 
              else if (local_pf_num == 0 && local_vf_num == 1376 && local_vf_active == 1) port_count[1376]++; 
              else if (local_pf_num == 0 && local_vf_num == 1377 && local_vf_active == 1) port_count[1377]++; 
              else if (local_pf_num == 0 && local_vf_num == 1378 && local_vf_active == 1) port_count[1378]++; 
              else if (local_pf_num == 0 && local_vf_num == 1379 && local_vf_active == 1) port_count[1379]++; 
              else if (local_pf_num == 0 && local_vf_num == 1380 && local_vf_active == 1) port_count[1380]++; 
              else if (local_pf_num == 0 && local_vf_num == 1381 && local_vf_active == 1) port_count[1381]++; 
              else if (local_pf_num == 0 && local_vf_num == 1382 && local_vf_active == 1) port_count[1382]++; 
              else if (local_pf_num == 0 && local_vf_num == 1383 && local_vf_active == 1) port_count[1383]++; 
              else if (local_pf_num == 0 && local_vf_num == 1384 && local_vf_active == 1) port_count[1384]++; 
              else if (local_pf_num == 0 && local_vf_num == 1385 && local_vf_active == 1) port_count[1385]++; 
              else if (local_pf_num == 0 && local_vf_num == 1386 && local_vf_active == 1) port_count[1386]++; 
              else if (local_pf_num == 0 && local_vf_num == 1387 && local_vf_active == 1) port_count[1387]++; 
              else if (local_pf_num == 0 && local_vf_num == 1388 && local_vf_active == 1) port_count[1388]++; 
              else if (local_pf_num == 0 && local_vf_num == 1389 && local_vf_active == 1) port_count[1389]++; 
              else if (local_pf_num == 0 && local_vf_num == 1390 && local_vf_active == 1) port_count[1390]++; 
              else if (local_pf_num == 0 && local_vf_num == 1391 && local_vf_active == 1) port_count[1391]++; 
              else if (local_pf_num == 0 && local_vf_num == 1392 && local_vf_active == 1) port_count[1392]++; 
              else if (local_pf_num == 0 && local_vf_num == 1393 && local_vf_active == 1) port_count[1393]++; 
              else if (local_pf_num == 0 && local_vf_num == 1394 && local_vf_active == 1) port_count[1394]++; 
              else if (local_pf_num == 0 && local_vf_num == 1395 && local_vf_active == 1) port_count[1395]++; 
              else if (local_pf_num == 0 && local_vf_num == 1396 && local_vf_active == 1) port_count[1396]++; 
              else if (local_pf_num == 0 && local_vf_num == 1397 && local_vf_active == 1) port_count[1397]++; 
              else if (local_pf_num == 0 && local_vf_num == 1398 && local_vf_active == 1) port_count[1398]++; 
              else if (local_pf_num == 0 && local_vf_num == 1399 && local_vf_active == 1) port_count[1399]++; 
              else if (local_pf_num == 0 && local_vf_num == 1400 && local_vf_active == 1) port_count[1400]++; 
              else if (local_pf_num == 0 && local_vf_num == 1401 && local_vf_active == 1) port_count[1401]++; 
              else if (local_pf_num == 0 && local_vf_num == 1402 && local_vf_active == 1) port_count[1402]++; 
              else if (local_pf_num == 0 && local_vf_num == 1403 && local_vf_active == 1) port_count[1403]++; 
              else if (local_pf_num == 0 && local_vf_num == 1404 && local_vf_active == 1) port_count[1404]++; 
              else if (local_pf_num == 0 && local_vf_num == 1405 && local_vf_active == 1) port_count[1405]++; 
              else if (local_pf_num == 0 && local_vf_num == 1406 && local_vf_active == 1) port_count[1406]++; 
              else if (local_pf_num == 0 && local_vf_num == 1407 && local_vf_active == 1) port_count[1407]++; 
              else if (local_pf_num == 0 && local_vf_num == 1408 && local_vf_active == 1) port_count[1408]++; 
              else if (local_pf_num == 0 && local_vf_num == 1409 && local_vf_active == 1) port_count[1409]++; 
              else if (local_pf_num == 0 && local_vf_num == 1410 && local_vf_active == 1) port_count[1410]++; 
              else if (local_pf_num == 0 && local_vf_num == 1411 && local_vf_active == 1) port_count[1411]++; 
              else if (local_pf_num == 0 && local_vf_num == 1412 && local_vf_active == 1) port_count[1412]++; 
              else if (local_pf_num == 0 && local_vf_num == 1413 && local_vf_active == 1) port_count[1413]++; 
              else if (local_pf_num == 0 && local_vf_num == 1414 && local_vf_active == 1) port_count[1414]++; 
              else if (local_pf_num == 0 && local_vf_num == 1415 && local_vf_active == 1) port_count[1415]++; 
              else if (local_pf_num == 0 && local_vf_num == 1416 && local_vf_active == 1) port_count[1416]++; 
              else if (local_pf_num == 0 && local_vf_num == 1417 && local_vf_active == 1) port_count[1417]++; 
              else if (local_pf_num == 0 && local_vf_num == 1418 && local_vf_active == 1) port_count[1418]++; 
              else if (local_pf_num == 0 && local_vf_num == 1419 && local_vf_active == 1) port_count[1419]++; 
              else if (local_pf_num == 0 && local_vf_num == 1420 && local_vf_active == 1) port_count[1420]++; 
              else if (local_pf_num == 0 && local_vf_num == 1421 && local_vf_active == 1) port_count[1421]++; 
              else if (local_pf_num == 0 && local_vf_num == 1422 && local_vf_active == 1) port_count[1422]++; 
              else if (local_pf_num == 0 && local_vf_num == 1423 && local_vf_active == 1) port_count[1423]++; 
              else if (local_pf_num == 0 && local_vf_num == 1424 && local_vf_active == 1) port_count[1424]++; 
              else if (local_pf_num == 0 && local_vf_num == 1425 && local_vf_active == 1) port_count[1425]++; 
              else if (local_pf_num == 0 && local_vf_num == 1426 && local_vf_active == 1) port_count[1426]++; 
              else if (local_pf_num == 0 && local_vf_num == 1427 && local_vf_active == 1) port_count[1427]++; 
              else if (local_pf_num == 0 && local_vf_num == 1428 && local_vf_active == 1) port_count[1428]++; 
              else if (local_pf_num == 0 && local_vf_num == 1429 && local_vf_active == 1) port_count[1429]++; 
              else if (local_pf_num == 0 && local_vf_num == 1430 && local_vf_active == 1) port_count[1430]++; 
              else if (local_pf_num == 0 && local_vf_num == 1431 && local_vf_active == 1) port_count[1431]++; 
              else if (local_pf_num == 0 && local_vf_num == 1432 && local_vf_active == 1) port_count[1432]++; 
              else if (local_pf_num == 0 && local_vf_num == 1433 && local_vf_active == 1) port_count[1433]++; 
              else if (local_pf_num == 0 && local_vf_num == 1434 && local_vf_active == 1) port_count[1434]++; 
              else if (local_pf_num == 0 && local_vf_num == 1435 && local_vf_active == 1) port_count[1435]++; 
              else if (local_pf_num == 0 && local_vf_num == 1436 && local_vf_active == 1) port_count[1436]++; 
              else if (local_pf_num == 0 && local_vf_num == 1437 && local_vf_active == 1) port_count[1437]++; 
              else if (local_pf_num == 0 && local_vf_num == 1438 && local_vf_active == 1) port_count[1438]++; 
              else if (local_pf_num == 0 && local_vf_num == 1439 && local_vf_active == 1) port_count[1439]++; 
              else if (local_pf_num == 0 && local_vf_num == 1440 && local_vf_active == 1) port_count[1440]++; 
              else if (local_pf_num == 0 && local_vf_num == 1441 && local_vf_active == 1) port_count[1441]++; 
              else if (local_pf_num == 0 && local_vf_num == 1442 && local_vf_active == 1) port_count[1442]++; 
              else if (local_pf_num == 0 && local_vf_num == 1443 && local_vf_active == 1) port_count[1443]++; 
              else if (local_pf_num == 0 && local_vf_num == 1444 && local_vf_active == 1) port_count[1444]++; 
              else if (local_pf_num == 0 && local_vf_num == 1445 && local_vf_active == 1) port_count[1445]++; 
              else if (local_pf_num == 0 && local_vf_num == 1446 && local_vf_active == 1) port_count[1446]++; 
              else if (local_pf_num == 0 && local_vf_num == 1447 && local_vf_active == 1) port_count[1447]++; 
              else if (local_pf_num == 0 && local_vf_num == 1448 && local_vf_active == 1) port_count[1448]++; 
              else if (local_pf_num == 0 && local_vf_num == 1449 && local_vf_active == 1) port_count[1449]++; 
              else if (local_pf_num == 0 && local_vf_num == 1450 && local_vf_active == 1) port_count[1450]++; 
              else if (local_pf_num == 0 && local_vf_num == 1451 && local_vf_active == 1) port_count[1451]++; 
              else if (local_pf_num == 0 && local_vf_num == 1452 && local_vf_active == 1) port_count[1452]++; 
              else if (local_pf_num == 0 && local_vf_num == 1453 && local_vf_active == 1) port_count[1453]++; 
              else if (local_pf_num == 0 && local_vf_num == 1454 && local_vf_active == 1) port_count[1454]++; 
              else if (local_pf_num == 0 && local_vf_num == 1455 && local_vf_active == 1) port_count[1455]++; 
              else if (local_pf_num == 0 && local_vf_num == 1456 && local_vf_active == 1) port_count[1456]++; 
              else if (local_pf_num == 0 && local_vf_num == 1457 && local_vf_active == 1) port_count[1457]++; 
              else if (local_pf_num == 0 && local_vf_num == 1458 && local_vf_active == 1) port_count[1458]++; 
              else if (local_pf_num == 0 && local_vf_num == 1459 && local_vf_active == 1) port_count[1459]++; 
              else if (local_pf_num == 0 && local_vf_num == 1460 && local_vf_active == 1) port_count[1460]++; 
              else if (local_pf_num == 0 && local_vf_num == 1461 && local_vf_active == 1) port_count[1461]++; 
              else if (local_pf_num == 0 && local_vf_num == 1462 && local_vf_active == 1) port_count[1462]++; 
              else if (local_pf_num == 0 && local_vf_num == 1463 && local_vf_active == 1) port_count[1463]++; 
              else if (local_pf_num == 0 && local_vf_num == 1464 && local_vf_active == 1) port_count[1464]++; 
              else if (local_pf_num == 0 && local_vf_num == 1465 && local_vf_active == 1) port_count[1465]++; 
              else if (local_pf_num == 0 && local_vf_num == 1466 && local_vf_active == 1) port_count[1466]++; 
              else if (local_pf_num == 0 && local_vf_num == 1467 && local_vf_active == 1) port_count[1467]++; 
              else if (local_pf_num == 0 && local_vf_num == 1468 && local_vf_active == 1) port_count[1468]++; 
              else if (local_pf_num == 0 && local_vf_num == 1469 && local_vf_active == 1) port_count[1469]++; 
              else if (local_pf_num == 0 && local_vf_num == 1470 && local_vf_active == 1) port_count[1470]++; 
              else if (local_pf_num == 0 && local_vf_num == 1471 && local_vf_active == 1) port_count[1471]++; 
              else if (local_pf_num == 0 && local_vf_num == 1472 && local_vf_active == 1) port_count[1472]++; 
              else if (local_pf_num == 0 && local_vf_num == 1473 && local_vf_active == 1) port_count[1473]++; 
              else if (local_pf_num == 0 && local_vf_num == 1474 && local_vf_active == 1) port_count[1474]++; 
              else if (local_pf_num == 0 && local_vf_num == 1475 && local_vf_active == 1) port_count[1475]++; 
              else if (local_pf_num == 0 && local_vf_num == 1476 && local_vf_active == 1) port_count[1476]++; 
              else if (local_pf_num == 0 && local_vf_num == 1477 && local_vf_active == 1) port_count[1477]++; 
              else if (local_pf_num == 0 && local_vf_num == 1478 && local_vf_active == 1) port_count[1478]++; 
              else if (local_pf_num == 0 && local_vf_num == 1479 && local_vf_active == 1) port_count[1479]++; 
              else if (local_pf_num == 0 && local_vf_num == 1480 && local_vf_active == 1) port_count[1480]++; 
              else if (local_pf_num == 0 && local_vf_num == 1481 && local_vf_active == 1) port_count[1481]++; 
              else if (local_pf_num == 0 && local_vf_num == 1482 && local_vf_active == 1) port_count[1482]++; 
              else if (local_pf_num == 0 && local_vf_num == 1483 && local_vf_active == 1) port_count[1483]++; 
              else if (local_pf_num == 0 && local_vf_num == 1484 && local_vf_active == 1) port_count[1484]++; 
              else if (local_pf_num == 0 && local_vf_num == 1485 && local_vf_active == 1) port_count[1485]++; 
              else if (local_pf_num == 0 && local_vf_num == 1486 && local_vf_active == 1) port_count[1486]++; 
              else if (local_pf_num == 0 && local_vf_num == 1487 && local_vf_active == 1) port_count[1487]++; 
              else if (local_pf_num == 0 && local_vf_num == 1488 && local_vf_active == 1) port_count[1488]++; 
              else if (local_pf_num == 0 && local_vf_num == 1489 && local_vf_active == 1) port_count[1489]++; 
              else if (local_pf_num == 0 && local_vf_num == 1490 && local_vf_active == 1) port_count[1490]++; 
              else if (local_pf_num == 0 && local_vf_num == 1491 && local_vf_active == 1) port_count[1491]++; 
              else if (local_pf_num == 0 && local_vf_num == 1492 && local_vf_active == 1) port_count[1492]++; 
              else if (local_pf_num == 0 && local_vf_num == 1493 && local_vf_active == 1) port_count[1493]++; 
              else if (local_pf_num == 0 && local_vf_num == 1494 && local_vf_active == 1) port_count[1494]++; 
              else if (local_pf_num == 0 && local_vf_num == 1495 && local_vf_active == 1) port_count[1495]++; 
              else if (local_pf_num == 0 && local_vf_num == 1496 && local_vf_active == 1) port_count[1496]++; 
              else if (local_pf_num == 0 && local_vf_num == 1497 && local_vf_active == 1) port_count[1497]++; 
              else if (local_pf_num == 0 && local_vf_num == 1498 && local_vf_active == 1) port_count[1498]++; 
              else if (local_pf_num == 0 && local_vf_num == 1499 && local_vf_active == 1) port_count[1499]++; 
              else if (local_pf_num == 0 && local_vf_num == 1500 && local_vf_active == 1) port_count[1500]++; 
              else if (local_pf_num == 0 && local_vf_num == 1501 && local_vf_active == 1) port_count[1501]++; 
              else if (local_pf_num == 0 && local_vf_num == 1502 && local_vf_active == 1) port_count[1502]++; 
              else if (local_pf_num == 0 && local_vf_num == 1503 && local_vf_active == 1) port_count[1503]++; 
              else if (local_pf_num == 0 && local_vf_num == 1504 && local_vf_active == 1) port_count[1504]++; 
              else if (local_pf_num == 0 && local_vf_num == 1505 && local_vf_active == 1) port_count[1505]++; 
              else if (local_pf_num == 0 && local_vf_num == 1506 && local_vf_active == 1) port_count[1506]++; 
              else if (local_pf_num == 0 && local_vf_num == 1507 && local_vf_active == 1) port_count[1507]++; 
              else if (local_pf_num == 0 && local_vf_num == 1508 && local_vf_active == 1) port_count[1508]++; 
              else if (local_pf_num == 0 && local_vf_num == 1509 && local_vf_active == 1) port_count[1509]++; 
              else if (local_pf_num == 0 && local_vf_num == 1510 && local_vf_active == 1) port_count[1510]++; 
              else if (local_pf_num == 0 && local_vf_num == 1511 && local_vf_active == 1) port_count[1511]++; 
              else if (local_pf_num == 0 && local_vf_num == 1512 && local_vf_active == 1) port_count[1512]++; 
              else if (local_pf_num == 0 && local_vf_num == 1513 && local_vf_active == 1) port_count[1513]++; 
              else if (local_pf_num == 0 && local_vf_num == 1514 && local_vf_active == 1) port_count[1514]++; 
              else if (local_pf_num == 0 && local_vf_num == 1515 && local_vf_active == 1) port_count[1515]++; 
              else if (local_pf_num == 0 && local_vf_num == 1516 && local_vf_active == 1) port_count[1516]++; 
              else if (local_pf_num == 0 && local_vf_num == 1517 && local_vf_active == 1) port_count[1517]++; 
              else if (local_pf_num == 0 && local_vf_num == 1518 && local_vf_active == 1) port_count[1518]++; 
              else if (local_pf_num == 0 && local_vf_num == 1519 && local_vf_active == 1) port_count[1519]++; 
              else if (local_pf_num == 0 && local_vf_num == 1520 && local_vf_active == 1) port_count[1520]++; 
              else if (local_pf_num == 0 && local_vf_num == 1521 && local_vf_active == 1) port_count[1521]++; 
              else if (local_pf_num == 0 && local_vf_num == 1522 && local_vf_active == 1) port_count[1522]++; 
              else if (local_pf_num == 0 && local_vf_num == 1523 && local_vf_active == 1) port_count[1523]++; 
              else if (local_pf_num == 0 && local_vf_num == 1524 && local_vf_active == 1) port_count[1524]++; 
              else if (local_pf_num == 0 && local_vf_num == 1525 && local_vf_active == 1) port_count[1525]++; 
              else if (local_pf_num == 0 && local_vf_num == 1526 && local_vf_active == 1) port_count[1526]++; 
              else if (local_pf_num == 0 && local_vf_num == 1527 && local_vf_active == 1) port_count[1527]++; 
              else if (local_pf_num == 0 && local_vf_num == 1528 && local_vf_active == 1) port_count[1528]++; 
              else if (local_pf_num == 0 && local_vf_num == 1529 && local_vf_active == 1) port_count[1529]++; 
              else if (local_pf_num == 0 && local_vf_num == 1530 && local_vf_active == 1) port_count[1530]++; 
              else if (local_pf_num == 0 && local_vf_num == 1531 && local_vf_active == 1) port_count[1531]++; 
              else if (local_pf_num == 0 && local_vf_num == 1532 && local_vf_active == 1) port_count[1532]++; 
              else if (local_pf_num == 0 && local_vf_num == 1533 && local_vf_active == 1) port_count[1533]++; 
              else if (local_pf_num == 0 && local_vf_num == 1534 && local_vf_active == 1) port_count[1534]++; 
              else if (local_pf_num == 0 && local_vf_num == 1535 && local_vf_active == 1) port_count[1535]++; 
              else if (local_pf_num == 0 && local_vf_num == 1536 && local_vf_active == 1) port_count[1536]++; 
              else if (local_pf_num == 0 && local_vf_num == 1537 && local_vf_active == 1) port_count[1537]++; 
              else if (local_pf_num == 0 && local_vf_num == 1538 && local_vf_active == 1) port_count[1538]++; 
              else if (local_pf_num == 0 && local_vf_num == 1539 && local_vf_active == 1) port_count[1539]++; 
              else if (local_pf_num == 0 && local_vf_num == 1540 && local_vf_active == 1) port_count[1540]++; 
              else if (local_pf_num == 0 && local_vf_num == 1541 && local_vf_active == 1) port_count[1541]++; 
              else if (local_pf_num == 0 && local_vf_num == 1542 && local_vf_active == 1) port_count[1542]++; 
              else if (local_pf_num == 0 && local_vf_num == 1543 && local_vf_active == 1) port_count[1543]++; 
              else if (local_pf_num == 0 && local_vf_num == 1544 && local_vf_active == 1) port_count[1544]++; 
              else if (local_pf_num == 0 && local_vf_num == 1545 && local_vf_active == 1) port_count[1545]++; 
              else if (local_pf_num == 0 && local_vf_num == 1546 && local_vf_active == 1) port_count[1546]++; 
              else if (local_pf_num == 0 && local_vf_num == 1547 && local_vf_active == 1) port_count[1547]++; 
              else if (local_pf_num == 0 && local_vf_num == 1548 && local_vf_active == 1) port_count[1548]++; 
              else if (local_pf_num == 0 && local_vf_num == 1549 && local_vf_active == 1) port_count[1549]++; 
              else if (local_pf_num == 0 && local_vf_num == 1550 && local_vf_active == 1) port_count[1550]++; 
              else if (local_pf_num == 0 && local_vf_num == 1551 && local_vf_active == 1) port_count[1551]++; 
              else if (local_pf_num == 0 && local_vf_num == 1552 && local_vf_active == 1) port_count[1552]++; 
              else if (local_pf_num == 0 && local_vf_num == 1553 && local_vf_active == 1) port_count[1553]++; 
              else if (local_pf_num == 0 && local_vf_num == 1554 && local_vf_active == 1) port_count[1554]++; 
              else if (local_pf_num == 0 && local_vf_num == 1555 && local_vf_active == 1) port_count[1555]++; 
              else if (local_pf_num == 0 && local_vf_num == 1556 && local_vf_active == 1) port_count[1556]++; 
              else if (local_pf_num == 0 && local_vf_num == 1557 && local_vf_active == 1) port_count[1557]++; 
              else if (local_pf_num == 0 && local_vf_num == 1558 && local_vf_active == 1) port_count[1558]++; 
              else if (local_pf_num == 0 && local_vf_num == 1559 && local_vf_active == 1) port_count[1559]++; 
              else if (local_pf_num == 0 && local_vf_num == 1560 && local_vf_active == 1) port_count[1560]++; 
              else if (local_pf_num == 0 && local_vf_num == 1561 && local_vf_active == 1) port_count[1561]++; 
              else if (local_pf_num == 0 && local_vf_num == 1562 && local_vf_active == 1) port_count[1562]++; 
              else if (local_pf_num == 0 && local_vf_num == 1563 && local_vf_active == 1) port_count[1563]++; 
              else if (local_pf_num == 0 && local_vf_num == 1564 && local_vf_active == 1) port_count[1564]++; 
              else if (local_pf_num == 0 && local_vf_num == 1565 && local_vf_active == 1) port_count[1565]++; 
              else if (local_pf_num == 0 && local_vf_num == 1566 && local_vf_active == 1) port_count[1566]++; 
              else if (local_pf_num == 0 && local_vf_num == 1567 && local_vf_active == 1) port_count[1567]++; 
              else if (local_pf_num == 0 && local_vf_num == 1568 && local_vf_active == 1) port_count[1568]++; 
              else if (local_pf_num == 0 && local_vf_num == 1569 && local_vf_active == 1) port_count[1569]++; 
              else if (local_pf_num == 0 && local_vf_num == 1570 && local_vf_active == 1) port_count[1570]++; 
              else if (local_pf_num == 0 && local_vf_num == 1571 && local_vf_active == 1) port_count[1571]++; 
              else if (local_pf_num == 0 && local_vf_num == 1572 && local_vf_active == 1) port_count[1572]++; 
              else if (local_pf_num == 0 && local_vf_num == 1573 && local_vf_active == 1) port_count[1573]++; 
              else if (local_pf_num == 0 && local_vf_num == 1574 && local_vf_active == 1) port_count[1574]++; 
              else if (local_pf_num == 0 && local_vf_num == 1575 && local_vf_active == 1) port_count[1575]++; 
              else if (local_pf_num == 0 && local_vf_num == 1576 && local_vf_active == 1) port_count[1576]++; 
              else if (local_pf_num == 0 && local_vf_num == 1577 && local_vf_active == 1) port_count[1577]++; 
              else if (local_pf_num == 0 && local_vf_num == 1578 && local_vf_active == 1) port_count[1578]++; 
              else if (local_pf_num == 0 && local_vf_num == 1579 && local_vf_active == 1) port_count[1579]++; 
              else if (local_pf_num == 0 && local_vf_num == 1580 && local_vf_active == 1) port_count[1580]++; 
              else if (local_pf_num == 0 && local_vf_num == 1581 && local_vf_active == 1) port_count[1581]++; 
              else if (local_pf_num == 0 && local_vf_num == 1582 && local_vf_active == 1) port_count[1582]++; 
              else if (local_pf_num == 0 && local_vf_num == 1583 && local_vf_active == 1) port_count[1583]++; 
              else if (local_pf_num == 0 && local_vf_num == 1584 && local_vf_active == 1) port_count[1584]++; 
              else if (local_pf_num == 0 && local_vf_num == 1585 && local_vf_active == 1) port_count[1585]++; 
              else if (local_pf_num == 0 && local_vf_num == 1586 && local_vf_active == 1) port_count[1586]++; 
              else if (local_pf_num == 0 && local_vf_num == 1587 && local_vf_active == 1) port_count[1587]++; 
              else if (local_pf_num == 0 && local_vf_num == 1588 && local_vf_active == 1) port_count[1588]++; 
              else if (local_pf_num == 0 && local_vf_num == 1589 && local_vf_active == 1) port_count[1589]++; 
              else if (local_pf_num == 0 && local_vf_num == 1590 && local_vf_active == 1) port_count[1590]++; 
              else if (local_pf_num == 0 && local_vf_num == 1591 && local_vf_active == 1) port_count[1591]++; 
              else if (local_pf_num == 0 && local_vf_num == 1592 && local_vf_active == 1) port_count[1592]++; 
              else if (local_pf_num == 0 && local_vf_num == 1593 && local_vf_active == 1) port_count[1593]++; 
              else if (local_pf_num == 0 && local_vf_num == 1594 && local_vf_active == 1) port_count[1594]++; 
              else if (local_pf_num == 0 && local_vf_num == 1595 && local_vf_active == 1) port_count[1595]++; 
              else if (local_pf_num == 0 && local_vf_num == 1596 && local_vf_active == 1) port_count[1596]++; 
              else if (local_pf_num == 0 && local_vf_num == 1597 && local_vf_active == 1) port_count[1597]++; 
              else if (local_pf_num == 0 && local_vf_num == 1598 && local_vf_active == 1) port_count[1598]++; 
              else if (local_pf_num == 0 && local_vf_num == 1599 && local_vf_active == 1) port_count[1599]++; 
              else if (local_pf_num == 0 && local_vf_num == 1600 && local_vf_active == 1) port_count[1600]++; 
              else if (local_pf_num == 0 && local_vf_num == 1601 && local_vf_active == 1) port_count[1601]++; 
              else if (local_pf_num == 0 && local_vf_num == 1602 && local_vf_active == 1) port_count[1602]++; 
              else if (local_pf_num == 0 && local_vf_num == 1603 && local_vf_active == 1) port_count[1603]++; 
              else if (local_pf_num == 0 && local_vf_num == 1604 && local_vf_active == 1) port_count[1604]++; 
              else if (local_pf_num == 0 && local_vf_num == 1605 && local_vf_active == 1) port_count[1605]++; 
              else if (local_pf_num == 0 && local_vf_num == 1606 && local_vf_active == 1) port_count[1606]++; 
              else if (local_pf_num == 0 && local_vf_num == 1607 && local_vf_active == 1) port_count[1607]++; 
              else if (local_pf_num == 0 && local_vf_num == 1608 && local_vf_active == 1) port_count[1608]++; 
              else if (local_pf_num == 0 && local_vf_num == 1609 && local_vf_active == 1) port_count[1609]++; 
              else if (local_pf_num == 0 && local_vf_num == 1610 && local_vf_active == 1) port_count[1610]++; 
              else if (local_pf_num == 0 && local_vf_num == 1611 && local_vf_active == 1) port_count[1611]++; 
              else if (local_pf_num == 0 && local_vf_num == 1612 && local_vf_active == 1) port_count[1612]++; 
              else if (local_pf_num == 0 && local_vf_num == 1613 && local_vf_active == 1) port_count[1613]++; 
              else if (local_pf_num == 0 && local_vf_num == 1614 && local_vf_active == 1) port_count[1614]++; 
              else if (local_pf_num == 0 && local_vf_num == 1615 && local_vf_active == 1) port_count[1615]++; 
              else if (local_pf_num == 0 && local_vf_num == 1616 && local_vf_active == 1) port_count[1616]++; 
              else if (local_pf_num == 0 && local_vf_num == 1617 && local_vf_active == 1) port_count[1617]++; 
              else if (local_pf_num == 0 && local_vf_num == 1618 && local_vf_active == 1) port_count[1618]++; 
              else if (local_pf_num == 0 && local_vf_num == 1619 && local_vf_active == 1) port_count[1619]++; 
              else if (local_pf_num == 0 && local_vf_num == 1620 && local_vf_active == 1) port_count[1620]++; 
              else if (local_pf_num == 0 && local_vf_num == 1621 && local_vf_active == 1) port_count[1621]++; 
              else if (local_pf_num == 0 && local_vf_num == 1622 && local_vf_active == 1) port_count[1622]++; 
              else if (local_pf_num == 0 && local_vf_num == 1623 && local_vf_active == 1) port_count[1623]++; 
              else if (local_pf_num == 0 && local_vf_num == 1624 && local_vf_active == 1) port_count[1624]++; 
              else if (local_pf_num == 0 && local_vf_num == 1625 && local_vf_active == 1) port_count[1625]++; 
              else if (local_pf_num == 0 && local_vf_num == 1626 && local_vf_active == 1) port_count[1626]++; 
              else if (local_pf_num == 0 && local_vf_num == 1627 && local_vf_active == 1) port_count[1627]++; 
              else if (local_pf_num == 0 && local_vf_num == 1628 && local_vf_active == 1) port_count[1628]++; 
              else if (local_pf_num == 0 && local_vf_num == 1629 && local_vf_active == 1) port_count[1629]++; 
              else if (local_pf_num == 0 && local_vf_num == 1630 && local_vf_active == 1) port_count[1630]++; 
              else if (local_pf_num == 0 && local_vf_num == 1631 && local_vf_active == 1) port_count[1631]++; 
              else if (local_pf_num == 0 && local_vf_num == 1632 && local_vf_active == 1) port_count[1632]++; 
              else if (local_pf_num == 0 && local_vf_num == 1633 && local_vf_active == 1) port_count[1633]++; 
              else if (local_pf_num == 0 && local_vf_num == 1634 && local_vf_active == 1) port_count[1634]++; 
              else if (local_pf_num == 0 && local_vf_num == 1635 && local_vf_active == 1) port_count[1635]++; 
              else if (local_pf_num == 0 && local_vf_num == 1636 && local_vf_active == 1) port_count[1636]++; 
              else if (local_pf_num == 0 && local_vf_num == 1637 && local_vf_active == 1) port_count[1637]++; 
              else if (local_pf_num == 0 && local_vf_num == 1638 && local_vf_active == 1) port_count[1638]++; 
              else if (local_pf_num == 0 && local_vf_num == 1639 && local_vf_active == 1) port_count[1639]++; 
              else if (local_pf_num == 0 && local_vf_num == 1640 && local_vf_active == 1) port_count[1640]++; 
              else if (local_pf_num == 0 && local_vf_num == 1641 && local_vf_active == 1) port_count[1641]++; 
              else if (local_pf_num == 0 && local_vf_num == 1642 && local_vf_active == 1) port_count[1642]++; 
              else if (local_pf_num == 0 && local_vf_num == 1643 && local_vf_active == 1) port_count[1643]++; 
              else if (local_pf_num == 0 && local_vf_num == 1644 && local_vf_active == 1) port_count[1644]++; 
              else if (local_pf_num == 0 && local_vf_num == 1645 && local_vf_active == 1) port_count[1645]++; 
              else if (local_pf_num == 0 && local_vf_num == 1646 && local_vf_active == 1) port_count[1646]++; 
              else if (local_pf_num == 0 && local_vf_num == 1647 && local_vf_active == 1) port_count[1647]++; 
              else if (local_pf_num == 0 && local_vf_num == 1648 && local_vf_active == 1) port_count[1648]++; 
              else if (local_pf_num == 0 && local_vf_num == 1649 && local_vf_active == 1) port_count[1649]++; 
              else if (local_pf_num == 0 && local_vf_num == 1650 && local_vf_active == 1) port_count[1650]++; 
              else if (local_pf_num == 0 && local_vf_num == 1651 && local_vf_active == 1) port_count[1651]++; 
              else if (local_pf_num == 0 && local_vf_num == 1652 && local_vf_active == 1) port_count[1652]++; 
              else if (local_pf_num == 0 && local_vf_num == 1653 && local_vf_active == 1) port_count[1653]++; 
              else if (local_pf_num == 0 && local_vf_num == 1654 && local_vf_active == 1) port_count[1654]++; 
              else if (local_pf_num == 0 && local_vf_num == 1655 && local_vf_active == 1) port_count[1655]++; 
              else if (local_pf_num == 0 && local_vf_num == 1656 && local_vf_active == 1) port_count[1656]++; 
              else if (local_pf_num == 0 && local_vf_num == 1657 && local_vf_active == 1) port_count[1657]++; 
              else if (local_pf_num == 0 && local_vf_num == 1658 && local_vf_active == 1) port_count[1658]++; 
              else if (local_pf_num == 0 && local_vf_num == 1659 && local_vf_active == 1) port_count[1659]++; 
              else if (local_pf_num == 0 && local_vf_num == 1660 && local_vf_active == 1) port_count[1660]++; 
              else if (local_pf_num == 0 && local_vf_num == 1661 && local_vf_active == 1) port_count[1661]++; 
              else if (local_pf_num == 0 && local_vf_num == 1662 && local_vf_active == 1) port_count[1662]++; 
              else if (local_pf_num == 0 && local_vf_num == 1663 && local_vf_active == 1) port_count[1663]++; 
              else if (local_pf_num == 0 && local_vf_num == 1664 && local_vf_active == 1) port_count[1664]++; 
              else if (local_pf_num == 0 && local_vf_num == 1665 && local_vf_active == 1) port_count[1665]++; 
              else if (local_pf_num == 0 && local_vf_num == 1666 && local_vf_active == 1) port_count[1666]++; 
              else if (local_pf_num == 0 && local_vf_num == 1667 && local_vf_active == 1) port_count[1667]++; 
              else if (local_pf_num == 0 && local_vf_num == 1668 && local_vf_active == 1) port_count[1668]++; 
              else if (local_pf_num == 0 && local_vf_num == 1669 && local_vf_active == 1) port_count[1669]++; 
              else if (local_pf_num == 0 && local_vf_num == 1670 && local_vf_active == 1) port_count[1670]++; 
              else if (local_pf_num == 0 && local_vf_num == 1671 && local_vf_active == 1) port_count[1671]++; 
              else if (local_pf_num == 0 && local_vf_num == 1672 && local_vf_active == 1) port_count[1672]++; 
              else if (local_pf_num == 0 && local_vf_num == 1673 && local_vf_active == 1) port_count[1673]++; 
              else if (local_pf_num == 0 && local_vf_num == 1674 && local_vf_active == 1) port_count[1674]++; 
              else if (local_pf_num == 0 && local_vf_num == 1675 && local_vf_active == 1) port_count[1675]++; 
              else if (local_pf_num == 0 && local_vf_num == 1676 && local_vf_active == 1) port_count[1676]++; 
              else if (local_pf_num == 0 && local_vf_num == 1677 && local_vf_active == 1) port_count[1677]++; 
              else if (local_pf_num == 0 && local_vf_num == 1678 && local_vf_active == 1) port_count[1678]++; 
              else if (local_pf_num == 0 && local_vf_num == 1679 && local_vf_active == 1) port_count[1679]++; 
              else if (local_pf_num == 0 && local_vf_num == 1680 && local_vf_active == 1) port_count[1680]++; 
              else if (local_pf_num == 0 && local_vf_num == 1681 && local_vf_active == 1) port_count[1681]++; 
              else if (local_pf_num == 0 && local_vf_num == 1682 && local_vf_active == 1) port_count[1682]++; 
              else if (local_pf_num == 0 && local_vf_num == 1683 && local_vf_active == 1) port_count[1683]++; 
              else if (local_pf_num == 0 && local_vf_num == 1684 && local_vf_active == 1) port_count[1684]++; 
              else if (local_pf_num == 0 && local_vf_num == 1685 && local_vf_active == 1) port_count[1685]++; 
              else if (local_pf_num == 0 && local_vf_num == 1686 && local_vf_active == 1) port_count[1686]++; 
              else if (local_pf_num == 0 && local_vf_num == 1687 && local_vf_active == 1) port_count[1687]++; 
              else if (local_pf_num == 0 && local_vf_num == 1688 && local_vf_active == 1) port_count[1688]++; 
              else if (local_pf_num == 0 && local_vf_num == 1689 && local_vf_active == 1) port_count[1689]++; 
              else if (local_pf_num == 0 && local_vf_num == 1690 && local_vf_active == 1) port_count[1690]++; 
              else if (local_pf_num == 0 && local_vf_num == 1691 && local_vf_active == 1) port_count[1691]++; 
              else if (local_pf_num == 0 && local_vf_num == 1692 && local_vf_active == 1) port_count[1692]++; 
              else if (local_pf_num == 0 && local_vf_num == 1693 && local_vf_active == 1) port_count[1693]++; 
              else if (local_pf_num == 0 && local_vf_num == 1694 && local_vf_active == 1) port_count[1694]++; 
              else if (local_pf_num == 0 && local_vf_num == 1695 && local_vf_active == 1) port_count[1695]++; 
              else if (local_pf_num == 0 && local_vf_num == 1696 && local_vf_active == 1) port_count[1696]++; 
              else if (local_pf_num == 0 && local_vf_num == 1697 && local_vf_active == 1) port_count[1697]++; 
              else if (local_pf_num == 0 && local_vf_num == 1698 && local_vf_active == 1) port_count[1698]++; 
              else if (local_pf_num == 0 && local_vf_num == 1699 && local_vf_active == 1) port_count[1699]++; 
              else if (local_pf_num == 0 && local_vf_num == 1700 && local_vf_active == 1) port_count[1700]++; 
              else if (local_pf_num == 0 && local_vf_num == 1701 && local_vf_active == 1) port_count[1701]++; 
              else if (local_pf_num == 0 && local_vf_num == 1702 && local_vf_active == 1) port_count[1702]++; 
              else if (local_pf_num == 0 && local_vf_num == 1703 && local_vf_active == 1) port_count[1703]++; 
              else if (local_pf_num == 0 && local_vf_num == 1704 && local_vf_active == 1) port_count[1704]++; 
              else if (local_pf_num == 0 && local_vf_num == 1705 && local_vf_active == 1) port_count[1705]++; 
              else if (local_pf_num == 0 && local_vf_num == 1706 && local_vf_active == 1) port_count[1706]++; 
              else if (local_pf_num == 0 && local_vf_num == 1707 && local_vf_active == 1) port_count[1707]++; 
              else if (local_pf_num == 0 && local_vf_num == 1708 && local_vf_active == 1) port_count[1708]++; 
              else if (local_pf_num == 0 && local_vf_num == 1709 && local_vf_active == 1) port_count[1709]++; 
              else if (local_pf_num == 0 && local_vf_num == 1710 && local_vf_active == 1) port_count[1710]++; 
              else if (local_pf_num == 0 && local_vf_num == 1711 && local_vf_active == 1) port_count[1711]++; 
              else if (local_pf_num == 0 && local_vf_num == 1712 && local_vf_active == 1) port_count[1712]++; 
              else if (local_pf_num == 0 && local_vf_num == 1713 && local_vf_active == 1) port_count[1713]++; 
              else if (local_pf_num == 0 && local_vf_num == 1714 && local_vf_active == 1) port_count[1714]++; 
              else if (local_pf_num == 0 && local_vf_num == 1715 && local_vf_active == 1) port_count[1715]++; 
              else if (local_pf_num == 0 && local_vf_num == 1716 && local_vf_active == 1) port_count[1716]++; 
              else if (local_pf_num == 0 && local_vf_num == 1717 && local_vf_active == 1) port_count[1717]++; 
              else if (local_pf_num == 0 && local_vf_num == 1718 && local_vf_active == 1) port_count[1718]++; 
              else if (local_pf_num == 0 && local_vf_num == 1719 && local_vf_active == 1) port_count[1719]++; 
              else if (local_pf_num == 0 && local_vf_num == 1720 && local_vf_active == 1) port_count[1720]++; 
              else if (local_pf_num == 0 && local_vf_num == 1721 && local_vf_active == 1) port_count[1721]++; 
              else if (local_pf_num == 0 && local_vf_num == 1722 && local_vf_active == 1) port_count[1722]++; 
              else if (local_pf_num == 0 && local_vf_num == 1723 && local_vf_active == 1) port_count[1723]++; 
              else if (local_pf_num == 0 && local_vf_num == 1724 && local_vf_active == 1) port_count[1724]++; 
              else if (local_pf_num == 0 && local_vf_num == 1725 && local_vf_active == 1) port_count[1725]++; 
              else if (local_pf_num == 0 && local_vf_num == 1726 && local_vf_active == 1) port_count[1726]++; 
              else if (local_pf_num == 0 && local_vf_num == 1727 && local_vf_active == 1) port_count[1727]++; 
              else if (local_pf_num == 0 && local_vf_num == 1728 && local_vf_active == 1) port_count[1728]++; 
              else if (local_pf_num == 0 && local_vf_num == 1729 && local_vf_active == 1) port_count[1729]++; 
              else if (local_pf_num == 0 && local_vf_num == 1730 && local_vf_active == 1) port_count[1730]++; 
              else if (local_pf_num == 0 && local_vf_num == 1731 && local_vf_active == 1) port_count[1731]++; 
              else if (local_pf_num == 0 && local_vf_num == 1732 && local_vf_active == 1) port_count[1732]++; 
              else if (local_pf_num == 0 && local_vf_num == 1733 && local_vf_active == 1) port_count[1733]++; 
              else if (local_pf_num == 0 && local_vf_num == 1734 && local_vf_active == 1) port_count[1734]++; 
              else if (local_pf_num == 0 && local_vf_num == 1735 && local_vf_active == 1) port_count[1735]++; 
              else if (local_pf_num == 0 && local_vf_num == 1736 && local_vf_active == 1) port_count[1736]++; 
              else if (local_pf_num == 0 && local_vf_num == 1737 && local_vf_active == 1) port_count[1737]++; 
              else if (local_pf_num == 0 && local_vf_num == 1738 && local_vf_active == 1) port_count[1738]++; 
              else if (local_pf_num == 0 && local_vf_num == 1739 && local_vf_active == 1) port_count[1739]++; 
              else if (local_pf_num == 0 && local_vf_num == 1740 && local_vf_active == 1) port_count[1740]++; 
              else if (local_pf_num == 0 && local_vf_num == 1741 && local_vf_active == 1) port_count[1741]++; 
              else if (local_pf_num == 0 && local_vf_num == 1742 && local_vf_active == 1) port_count[1742]++; 
              else if (local_pf_num == 0 && local_vf_num == 1743 && local_vf_active == 1) port_count[1743]++; 
              else if (local_pf_num == 0 && local_vf_num == 1744 && local_vf_active == 1) port_count[1744]++; 
              else if (local_pf_num == 0 && local_vf_num == 1745 && local_vf_active == 1) port_count[1745]++; 
              else if (local_pf_num == 0 && local_vf_num == 1746 && local_vf_active == 1) port_count[1746]++; 
              else if (local_pf_num == 0 && local_vf_num == 1747 && local_vf_active == 1) port_count[1747]++; 
              else if (local_pf_num == 0 && local_vf_num == 1748 && local_vf_active == 1) port_count[1748]++; 
              else if (local_pf_num == 0 && local_vf_num == 1749 && local_vf_active == 1) port_count[1749]++; 
              else if (local_pf_num == 0 && local_vf_num == 1750 && local_vf_active == 1) port_count[1750]++; 
              else if (local_pf_num == 0 && local_vf_num == 1751 && local_vf_active == 1) port_count[1751]++; 
              else if (local_pf_num == 0 && local_vf_num == 1752 && local_vf_active == 1) port_count[1752]++; 
              else if (local_pf_num == 0 && local_vf_num == 1753 && local_vf_active == 1) port_count[1753]++; 
              else if (local_pf_num == 0 && local_vf_num == 1754 && local_vf_active == 1) port_count[1754]++; 
              else if (local_pf_num == 0 && local_vf_num == 1755 && local_vf_active == 1) port_count[1755]++; 
              else if (local_pf_num == 0 && local_vf_num == 1756 && local_vf_active == 1) port_count[1756]++; 
              else if (local_pf_num == 0 && local_vf_num == 1757 && local_vf_active == 1) port_count[1757]++; 
              else if (local_pf_num == 0 && local_vf_num == 1758 && local_vf_active == 1) port_count[1758]++; 
              else if (local_pf_num == 0 && local_vf_num == 1759 && local_vf_active == 1) port_count[1759]++; 
              else if (local_pf_num == 0 && local_vf_num == 1760 && local_vf_active == 1) port_count[1760]++; 
              else if (local_pf_num == 0 && local_vf_num == 1761 && local_vf_active == 1) port_count[1761]++; 
              else if (local_pf_num == 0 && local_vf_num == 1762 && local_vf_active == 1) port_count[1762]++; 
              else if (local_pf_num == 0 && local_vf_num == 1763 && local_vf_active == 1) port_count[1763]++; 
              else if (local_pf_num == 0 && local_vf_num == 1764 && local_vf_active == 1) port_count[1764]++; 
              else if (local_pf_num == 0 && local_vf_num == 1765 && local_vf_active == 1) port_count[1765]++; 
              else if (local_pf_num == 0 && local_vf_num == 1766 && local_vf_active == 1) port_count[1766]++; 
              else if (local_pf_num == 0 && local_vf_num == 1767 && local_vf_active == 1) port_count[1767]++; 
              else if (local_pf_num == 0 && local_vf_num == 1768 && local_vf_active == 1) port_count[1768]++; 
              else if (local_pf_num == 0 && local_vf_num == 1769 && local_vf_active == 1) port_count[1769]++; 
              else if (local_pf_num == 0 && local_vf_num == 1770 && local_vf_active == 1) port_count[1770]++; 
              else if (local_pf_num == 0 && local_vf_num == 1771 && local_vf_active == 1) port_count[1771]++; 
              else if (local_pf_num == 0 && local_vf_num == 1772 && local_vf_active == 1) port_count[1772]++; 
              else if (local_pf_num == 0 && local_vf_num == 1773 && local_vf_active == 1) port_count[1773]++; 
              else if (local_pf_num == 0 && local_vf_num == 1774 && local_vf_active == 1) port_count[1774]++; 
              else if (local_pf_num == 0 && local_vf_num == 1775 && local_vf_active == 1) port_count[1775]++; 
              else if (local_pf_num == 0 && local_vf_num == 1776 && local_vf_active == 1) port_count[1776]++; 
              else if (local_pf_num == 0 && local_vf_num == 1777 && local_vf_active == 1) port_count[1777]++; 
              else if (local_pf_num == 0 && local_vf_num == 1778 && local_vf_active == 1) port_count[1778]++; 
              else if (local_pf_num == 0 && local_vf_num == 1779 && local_vf_active == 1) port_count[1779]++; 
              else if (local_pf_num == 0 && local_vf_num == 1780 && local_vf_active == 1) port_count[1780]++; 
              else if (local_pf_num == 0 && local_vf_num == 1781 && local_vf_active == 1) port_count[1781]++; 
              else if (local_pf_num == 0 && local_vf_num == 1782 && local_vf_active == 1) port_count[1782]++; 
              else if (local_pf_num == 0 && local_vf_num == 1783 && local_vf_active == 1) port_count[1783]++; 
              else if (local_pf_num == 0 && local_vf_num == 1784 && local_vf_active == 1) port_count[1784]++; 
              else if (local_pf_num == 0 && local_vf_num == 1785 && local_vf_active == 1) port_count[1785]++; 
              else if (local_pf_num == 0 && local_vf_num == 1786 && local_vf_active == 1) port_count[1786]++; 
              else if (local_pf_num == 0 && local_vf_num == 1787 && local_vf_active == 1) port_count[1787]++; 
              else if (local_pf_num == 0 && local_vf_num == 1788 && local_vf_active == 1) port_count[1788]++; 
              else if (local_pf_num == 0 && local_vf_num == 1789 && local_vf_active == 1) port_count[1789]++; 
              else if (local_pf_num == 0 && local_vf_num == 1790 && local_vf_active == 1) port_count[1790]++; 
              else if (local_pf_num == 0 && local_vf_num == 1791 && local_vf_active == 1) port_count[1791]++; 
              else if (local_pf_num == 0 && local_vf_num == 1792 && local_vf_active == 1) port_count[1792]++; 
              else if (local_pf_num == 0 && local_vf_num == 1793 && local_vf_active == 1) port_count[1793]++; 
              else if (local_pf_num == 0 && local_vf_num == 1794 && local_vf_active == 1) port_count[1794]++; 
              else if (local_pf_num == 0 && local_vf_num == 1795 && local_vf_active == 1) port_count[1795]++; 
              else if (local_pf_num == 0 && local_vf_num == 1796 && local_vf_active == 1) port_count[1796]++; 
              else if (local_pf_num == 0 && local_vf_num == 1797 && local_vf_active == 1) port_count[1797]++; 
              else if (local_pf_num == 0 && local_vf_num == 1798 && local_vf_active == 1) port_count[1798]++; 
              else if (local_pf_num == 0 && local_vf_num == 1799 && local_vf_active == 1) port_count[1799]++; 
              else if (local_pf_num == 0 && local_vf_num == 1800 && local_vf_active == 1) port_count[1800]++; 
              else if (local_pf_num == 0 && local_vf_num == 1801 && local_vf_active == 1) port_count[1801]++; 
              else if (local_pf_num == 0 && local_vf_num == 1802 && local_vf_active == 1) port_count[1802]++; 
              else if (local_pf_num == 0 && local_vf_num == 1803 && local_vf_active == 1) port_count[1803]++; 
              else if (local_pf_num == 0 && local_vf_num == 1804 && local_vf_active == 1) port_count[1804]++; 
              else if (local_pf_num == 0 && local_vf_num == 1805 && local_vf_active == 1) port_count[1805]++; 
              else if (local_pf_num == 0 && local_vf_num == 1806 && local_vf_active == 1) port_count[1806]++; 
              else if (local_pf_num == 0 && local_vf_num == 1807 && local_vf_active == 1) port_count[1807]++; 
              else if (local_pf_num == 0 && local_vf_num == 1808 && local_vf_active == 1) port_count[1808]++; 
              else if (local_pf_num == 0 && local_vf_num == 1809 && local_vf_active == 1) port_count[1809]++; 
              else if (local_pf_num == 0 && local_vf_num == 1810 && local_vf_active == 1) port_count[1810]++; 
              else if (local_pf_num == 0 && local_vf_num == 1811 && local_vf_active == 1) port_count[1811]++; 
              else if (local_pf_num == 0 && local_vf_num == 1812 && local_vf_active == 1) port_count[1812]++; 
              else if (local_pf_num == 0 && local_vf_num == 1813 && local_vf_active == 1) port_count[1813]++; 
              else if (local_pf_num == 0 && local_vf_num == 1814 && local_vf_active == 1) port_count[1814]++; 
              else if (local_pf_num == 0 && local_vf_num == 1815 && local_vf_active == 1) port_count[1815]++; 
              else if (local_pf_num == 0 && local_vf_num == 1816 && local_vf_active == 1) port_count[1816]++; 
              else if (local_pf_num == 0 && local_vf_num == 1817 && local_vf_active == 1) port_count[1817]++; 
              else if (local_pf_num == 0 && local_vf_num == 1818 && local_vf_active == 1) port_count[1818]++; 
              else if (local_pf_num == 0 && local_vf_num == 1819 && local_vf_active == 1) port_count[1819]++; 
              else if (local_pf_num == 0 && local_vf_num == 1820 && local_vf_active == 1) port_count[1820]++; 
              else if (local_pf_num == 0 && local_vf_num == 1821 && local_vf_active == 1) port_count[1821]++; 
              else if (local_pf_num == 0 && local_vf_num == 1822 && local_vf_active == 1) port_count[1822]++; 
              else if (local_pf_num == 0 && local_vf_num == 1823 && local_vf_active == 1) port_count[1823]++; 
              else if (local_pf_num == 0 && local_vf_num == 1824 && local_vf_active == 1) port_count[1824]++; 
              else if (local_pf_num == 0 && local_vf_num == 1825 && local_vf_active == 1) port_count[1825]++; 
              else if (local_pf_num == 0 && local_vf_num == 1826 && local_vf_active == 1) port_count[1826]++; 
              else if (local_pf_num == 0 && local_vf_num == 1827 && local_vf_active == 1) port_count[1827]++; 
              else if (local_pf_num == 0 && local_vf_num == 1828 && local_vf_active == 1) port_count[1828]++; 
              else if (local_pf_num == 0 && local_vf_num == 1829 && local_vf_active == 1) port_count[1829]++; 
              else if (local_pf_num == 0 && local_vf_num == 1830 && local_vf_active == 1) port_count[1830]++; 
              else if (local_pf_num == 0 && local_vf_num == 1831 && local_vf_active == 1) port_count[1831]++; 
              else if (local_pf_num == 0 && local_vf_num == 1832 && local_vf_active == 1) port_count[1832]++; 
              else if (local_pf_num == 0 && local_vf_num == 1833 && local_vf_active == 1) port_count[1833]++; 
              else if (local_pf_num == 0 && local_vf_num == 1834 && local_vf_active == 1) port_count[1834]++; 
              else if (local_pf_num == 0 && local_vf_num == 1835 && local_vf_active == 1) port_count[1835]++; 
              else if (local_pf_num == 0 && local_vf_num == 1836 && local_vf_active == 1) port_count[1836]++; 
              else if (local_pf_num == 0 && local_vf_num == 1837 && local_vf_active == 1) port_count[1837]++; 
              else if (local_pf_num == 0 && local_vf_num == 1838 && local_vf_active == 1) port_count[1838]++; 
              else if (local_pf_num == 0 && local_vf_num == 1839 && local_vf_active == 1) port_count[1839]++; 
              else if (local_pf_num == 0 && local_vf_num == 1840 && local_vf_active == 1) port_count[1840]++; 
              else if (local_pf_num == 0 && local_vf_num == 1841 && local_vf_active == 1) port_count[1841]++; 
              else if (local_pf_num == 0 && local_vf_num == 1842 && local_vf_active == 1) port_count[1842]++; 
              else if (local_pf_num == 0 && local_vf_num == 1843 && local_vf_active == 1) port_count[1843]++; 
              else if (local_pf_num == 0 && local_vf_num == 1844 && local_vf_active == 1) port_count[1844]++; 
              else if (local_pf_num == 0 && local_vf_num == 1845 && local_vf_active == 1) port_count[1845]++; 
              else if (local_pf_num == 0 && local_vf_num == 1846 && local_vf_active == 1) port_count[1846]++; 
              else if (local_pf_num == 0 && local_vf_num == 1847 && local_vf_active == 1) port_count[1847]++; 
              else if (local_pf_num == 0 && local_vf_num == 1848 && local_vf_active == 1) port_count[1848]++; 
              else if (local_pf_num == 0 && local_vf_num == 1849 && local_vf_active == 1) port_count[1849]++; 
              else if (local_pf_num == 0 && local_vf_num == 1850 && local_vf_active == 1) port_count[1850]++; 
              else if (local_pf_num == 0 && local_vf_num == 1851 && local_vf_active == 1) port_count[1851]++; 
              else if (local_pf_num == 0 && local_vf_num == 1852 && local_vf_active == 1) port_count[1852]++; 
              else if (local_pf_num == 0 && local_vf_num == 1853 && local_vf_active == 1) port_count[1853]++; 
              else if (local_pf_num == 0 && local_vf_num == 1854 && local_vf_active == 1) port_count[1854]++; 
              else if (local_pf_num == 0 && local_vf_num == 1855 && local_vf_active == 1) port_count[1855]++; 
              else if (local_pf_num == 0 && local_vf_num == 1856 && local_vf_active == 1) port_count[1856]++; 
              else if (local_pf_num == 0 && local_vf_num == 1857 && local_vf_active == 1) port_count[1857]++; 
              else if (local_pf_num == 0 && local_vf_num == 1858 && local_vf_active == 1) port_count[1858]++; 
              else if (local_pf_num == 0 && local_vf_num == 1859 && local_vf_active == 1) port_count[1859]++; 
              else if (local_pf_num == 0 && local_vf_num == 1860 && local_vf_active == 1) port_count[1860]++; 
              else if (local_pf_num == 0 && local_vf_num == 1861 && local_vf_active == 1) port_count[1861]++; 
              else if (local_pf_num == 0 && local_vf_num == 1862 && local_vf_active == 1) port_count[1862]++; 
              else if (local_pf_num == 0 && local_vf_num == 1863 && local_vf_active == 1) port_count[1863]++; 
              else if (local_pf_num == 0 && local_vf_num == 1864 && local_vf_active == 1) port_count[1864]++; 
              else if (local_pf_num == 0 && local_vf_num == 1865 && local_vf_active == 1) port_count[1865]++; 
              else if (local_pf_num == 0 && local_vf_num == 1866 && local_vf_active == 1) port_count[1866]++; 
              else if (local_pf_num == 0 && local_vf_num == 1867 && local_vf_active == 1) port_count[1867]++; 
              else if (local_pf_num == 0 && local_vf_num == 1868 && local_vf_active == 1) port_count[1868]++; 
              else if (local_pf_num == 0 && local_vf_num == 1869 && local_vf_active == 1) port_count[1869]++; 
              else if (local_pf_num == 0 && local_vf_num == 1870 && local_vf_active == 1) port_count[1870]++; 
              else if (local_pf_num == 0 && local_vf_num == 1871 && local_vf_active == 1) port_count[1871]++; 
              else if (local_pf_num == 0 && local_vf_num == 1872 && local_vf_active == 1) port_count[1872]++; 
              else if (local_pf_num == 0 && local_vf_num == 1873 && local_vf_active == 1) port_count[1873]++; 
              else if (local_pf_num == 0 && local_vf_num == 1874 && local_vf_active == 1) port_count[1874]++; 
              else if (local_pf_num == 0 && local_vf_num == 1875 && local_vf_active == 1) port_count[1875]++; 
              else if (local_pf_num == 0 && local_vf_num == 1876 && local_vf_active == 1) port_count[1876]++; 
              else if (local_pf_num == 0 && local_vf_num == 1877 && local_vf_active == 1) port_count[1877]++; 
              else if (local_pf_num == 0 && local_vf_num == 1878 && local_vf_active == 1) port_count[1878]++; 
              else if (local_pf_num == 0 && local_vf_num == 1879 && local_vf_active == 1) port_count[1879]++; 
              else if (local_pf_num == 0 && local_vf_num == 1880 && local_vf_active == 1) port_count[1880]++; 
              else if (local_pf_num == 0 && local_vf_num == 1881 && local_vf_active == 1) port_count[1881]++; 
              else if (local_pf_num == 0 && local_vf_num == 1882 && local_vf_active == 1) port_count[1882]++; 
              else if (local_pf_num == 0 && local_vf_num == 1883 && local_vf_active == 1) port_count[1883]++; 
              else if (local_pf_num == 0 && local_vf_num == 1884 && local_vf_active == 1) port_count[1884]++; 
              else if (local_pf_num == 0 && local_vf_num == 1885 && local_vf_active == 1) port_count[1885]++; 
              else if (local_pf_num == 0 && local_vf_num == 1886 && local_vf_active == 1) port_count[1886]++; 
              else if (local_pf_num == 0 && local_vf_num == 1887 && local_vf_active == 1) port_count[1887]++; 
              else if (local_pf_num == 0 && local_vf_num == 1888 && local_vf_active == 1) port_count[1888]++; 
              else if (local_pf_num == 0 && local_vf_num == 1889 && local_vf_active == 1) port_count[1889]++; 
              else if (local_pf_num == 0 && local_vf_num == 1890 && local_vf_active == 1) port_count[1890]++; 
              else if (local_pf_num == 0 && local_vf_num == 1891 && local_vf_active == 1) port_count[1891]++; 
              else if (local_pf_num == 0 && local_vf_num == 1892 && local_vf_active == 1) port_count[1892]++; 
              else if (local_pf_num == 0 && local_vf_num == 1893 && local_vf_active == 1) port_count[1893]++; 
              else if (local_pf_num == 0 && local_vf_num == 1894 && local_vf_active == 1) port_count[1894]++; 
              else if (local_pf_num == 0 && local_vf_num == 1895 && local_vf_active == 1) port_count[1895]++; 
              else if (local_pf_num == 0 && local_vf_num == 1896 && local_vf_active == 1) port_count[1896]++; 
              else if (local_pf_num == 0 && local_vf_num == 1897 && local_vf_active == 1) port_count[1897]++; 
              else if (local_pf_num == 0 && local_vf_num == 1898 && local_vf_active == 1) port_count[1898]++; 
              else if (local_pf_num == 0 && local_vf_num == 1899 && local_vf_active == 1) port_count[1899]++; 
              else if (local_pf_num == 0 && local_vf_num == 1900 && local_vf_active == 1) port_count[1900]++; 
              else if (local_pf_num == 0 && local_vf_num == 1901 && local_vf_active == 1) port_count[1901]++; 
              else if (local_pf_num == 0 && local_vf_num == 1902 && local_vf_active == 1) port_count[1902]++; 
              else if (local_pf_num == 0 && local_vf_num == 1903 && local_vf_active == 1) port_count[1903]++; 
              else if (local_pf_num == 0 && local_vf_num == 1904 && local_vf_active == 1) port_count[1904]++; 
              else if (local_pf_num == 0 && local_vf_num == 1905 && local_vf_active == 1) port_count[1905]++; 
              else if (local_pf_num == 0 && local_vf_num == 1906 && local_vf_active == 1) port_count[1906]++; 
              else if (local_pf_num == 0 && local_vf_num == 1907 && local_vf_active == 1) port_count[1907]++; 
              else if (local_pf_num == 0 && local_vf_num == 1908 && local_vf_active == 1) port_count[1908]++; 
              else if (local_pf_num == 0 && local_vf_num == 1909 && local_vf_active == 1) port_count[1909]++; 
              else if (local_pf_num == 0 && local_vf_num == 1910 && local_vf_active == 1) port_count[1910]++; 
              else if (local_pf_num == 0 && local_vf_num == 1911 && local_vf_active == 1) port_count[1911]++; 
              else if (local_pf_num == 0 && local_vf_num == 1912 && local_vf_active == 1) port_count[1912]++; 
              else if (local_pf_num == 0 && local_vf_num == 1913 && local_vf_active == 1) port_count[1913]++; 
              else if (local_pf_num == 0 && local_vf_num == 1914 && local_vf_active == 1) port_count[1914]++; 
              else if (local_pf_num == 0 && local_vf_num == 1915 && local_vf_active == 1) port_count[1915]++; 
              else if (local_pf_num == 0 && local_vf_num == 1916 && local_vf_active == 1) port_count[1916]++; 
              else if (local_pf_num == 0 && local_vf_num == 1917 && local_vf_active == 1) port_count[1917]++; 
              else if (local_pf_num == 0 && local_vf_num == 1918 && local_vf_active == 1) port_count[1918]++; 
              else if (local_pf_num == 0 && local_vf_num == 1919 && local_vf_active == 1) port_count[1919]++; 
              else if (local_pf_num == 0 && local_vf_num == 1920 && local_vf_active == 1) port_count[1920]++; 
              else if (local_pf_num == 0 && local_vf_num == 1921 && local_vf_active == 1) port_count[1921]++; 
              else if (local_pf_num == 0 && local_vf_num == 1922 && local_vf_active == 1) port_count[1922]++; 
              else if (local_pf_num == 0 && local_vf_num == 1923 && local_vf_active == 1) port_count[1923]++; 
              else if (local_pf_num == 0 && local_vf_num == 1924 && local_vf_active == 1) port_count[1924]++; 
              else if (local_pf_num == 0 && local_vf_num == 1925 && local_vf_active == 1) port_count[1925]++; 
              else if (local_pf_num == 0 && local_vf_num == 1926 && local_vf_active == 1) port_count[1926]++; 
              else if (local_pf_num == 0 && local_vf_num == 1927 && local_vf_active == 1) port_count[1927]++; 
              else if (local_pf_num == 0 && local_vf_num == 1928 && local_vf_active == 1) port_count[1928]++; 
              else if (local_pf_num == 0 && local_vf_num == 1929 && local_vf_active == 1) port_count[1929]++; 
              else if (local_pf_num == 0 && local_vf_num == 1930 && local_vf_active == 1) port_count[1930]++; 
              else if (local_pf_num == 0 && local_vf_num == 1931 && local_vf_active == 1) port_count[1931]++; 
              else if (local_pf_num == 0 && local_vf_num == 1932 && local_vf_active == 1) port_count[1932]++; 
              else if (local_pf_num == 0 && local_vf_num == 1933 && local_vf_active == 1) port_count[1933]++; 
              else if (local_pf_num == 0 && local_vf_num == 1934 && local_vf_active == 1) port_count[1934]++; 
              else if (local_pf_num == 0 && local_vf_num == 1935 && local_vf_active == 1) port_count[1935]++; 
              else if (local_pf_num == 0 && local_vf_num == 1936 && local_vf_active == 1) port_count[1936]++; 
              else if (local_pf_num == 0 && local_vf_num == 1937 && local_vf_active == 1) port_count[1937]++; 
              else if (local_pf_num == 0 && local_vf_num == 1938 && local_vf_active == 1) port_count[1938]++; 
              else if (local_pf_num == 0 && local_vf_num == 1939 && local_vf_active == 1) port_count[1939]++; 
              else if (local_pf_num == 0 && local_vf_num == 1940 && local_vf_active == 1) port_count[1940]++; 
              else if (local_pf_num == 0 && local_vf_num == 1941 && local_vf_active == 1) port_count[1941]++; 
              else if (local_pf_num == 0 && local_vf_num == 1942 && local_vf_active == 1) port_count[1942]++; 
              else if (local_pf_num == 0 && local_vf_num == 1943 && local_vf_active == 1) port_count[1943]++; 
              else if (local_pf_num == 0 && local_vf_num == 1944 && local_vf_active == 1) port_count[1944]++; 
              else if (local_pf_num == 0 && local_vf_num == 1945 && local_vf_active == 1) port_count[1945]++; 
              else if (local_pf_num == 0 && local_vf_num == 1946 && local_vf_active == 1) port_count[1946]++; 
              else if (local_pf_num == 0 && local_vf_num == 1947 && local_vf_active == 1) port_count[1947]++; 
              else if (local_pf_num == 0 && local_vf_num == 1948 && local_vf_active == 1) port_count[1948]++; 
              else if (local_pf_num == 0 && local_vf_num == 1949 && local_vf_active == 1) port_count[1949]++; 
              else if (local_pf_num == 0 && local_vf_num == 1950 && local_vf_active == 1) port_count[1950]++; 
              else if (local_pf_num == 0 && local_vf_num == 1951 && local_vf_active == 1) port_count[1951]++; 
              else if (local_pf_num == 0 && local_vf_num == 1952 && local_vf_active == 1) port_count[1952]++; 
              else if (local_pf_num == 0 && local_vf_num == 1953 && local_vf_active == 1) port_count[1953]++; 
              else if (local_pf_num == 0 && local_vf_num == 1954 && local_vf_active == 1) port_count[1954]++; 
              else if (local_pf_num == 0 && local_vf_num == 1955 && local_vf_active == 1) port_count[1955]++; 
              else if (local_pf_num == 0 && local_vf_num == 1956 && local_vf_active == 1) port_count[1956]++; 
              else if (local_pf_num == 0 && local_vf_num == 1957 && local_vf_active == 1) port_count[1957]++; 
              else if (local_pf_num == 0 && local_vf_num == 1958 && local_vf_active == 1) port_count[1958]++; 
              else if (local_pf_num == 0 && local_vf_num == 1959 && local_vf_active == 1) port_count[1959]++; 
              else if (local_pf_num == 0 && local_vf_num == 1960 && local_vf_active == 1) port_count[1960]++; 
              else if (local_pf_num == 0 && local_vf_num == 1961 && local_vf_active == 1) port_count[1961]++; 
              else if (local_pf_num == 0 && local_vf_num == 1962 && local_vf_active == 1) port_count[1962]++; 
              else if (local_pf_num == 0 && local_vf_num == 1963 && local_vf_active == 1) port_count[1963]++; 
              else if (local_pf_num == 0 && local_vf_num == 1964 && local_vf_active == 1) port_count[1964]++; 
              else if (local_pf_num == 0 && local_vf_num == 1965 && local_vf_active == 1) port_count[1965]++; 
              else if (local_pf_num == 0 && local_vf_num == 1966 && local_vf_active == 1) port_count[1966]++; 
              else if (local_pf_num == 0 && local_vf_num == 1967 && local_vf_active == 1) port_count[1967]++; 
              else if (local_pf_num == 0 && local_vf_num == 1968 && local_vf_active == 1) port_count[1968]++; 
              else if (local_pf_num == 0 && local_vf_num == 1969 && local_vf_active == 1) port_count[1969]++; 
              else if (local_pf_num == 0 && local_vf_num == 1970 && local_vf_active == 1) port_count[1970]++; 
              else if (local_pf_num == 0 && local_vf_num == 1971 && local_vf_active == 1) port_count[1971]++; 
              else if (local_pf_num == 0 && local_vf_num == 1972 && local_vf_active == 1) port_count[1972]++; 
              else if (local_pf_num == 0 && local_vf_num == 1973 && local_vf_active == 1) port_count[1973]++; 
              else if (local_pf_num == 0 && local_vf_num == 1974 && local_vf_active == 1) port_count[1974]++; 
              else if (local_pf_num == 0 && local_vf_num == 1975 && local_vf_active == 1) port_count[1975]++; 
              else if (local_pf_num == 0 && local_vf_num == 1976 && local_vf_active == 1) port_count[1976]++; 
              else if (local_pf_num == 0 && local_vf_num == 1977 && local_vf_active == 1) port_count[1977]++; 
              else if (local_pf_num == 0 && local_vf_num == 1978 && local_vf_active == 1) port_count[1978]++; 
              else if (local_pf_num == 0 && local_vf_num == 1979 && local_vf_active == 1) port_count[1979]++; 
              else if (local_pf_num == 0 && local_vf_num == 1980 && local_vf_active == 1) port_count[1980]++; 
              else if (local_pf_num == 0 && local_vf_num == 1981 && local_vf_active == 1) port_count[1981]++; 
              else if (local_pf_num == 0 && local_vf_num == 1982 && local_vf_active == 1) port_count[1982]++; 
              else if (local_pf_num == 0 && local_vf_num == 1983 && local_vf_active == 1) port_count[1983]++; 
              else if (local_pf_num == 0 && local_vf_num == 1984 && local_vf_active == 1) port_count[1984]++; 
              else if (local_pf_num == 0 && local_vf_num == 1985 && local_vf_active == 1) port_count[1985]++; 
              else if (local_pf_num == 0 && local_vf_num == 1986 && local_vf_active == 1) port_count[1986]++; 
              else if (local_pf_num == 0 && local_vf_num == 1987 && local_vf_active == 1) port_count[1987]++; 
              else if (local_pf_num == 0 && local_vf_num == 1988 && local_vf_active == 1) port_count[1988]++; 
              else if (local_pf_num == 0 && local_vf_num == 1989 && local_vf_active == 1) port_count[1989]++; 
              else if (local_pf_num == 0 && local_vf_num == 1990 && local_vf_active == 1) port_count[1990]++; 
              else if (local_pf_num == 0 && local_vf_num == 1991 && local_vf_active == 1) port_count[1991]++; 
              else if (local_pf_num == 0 && local_vf_num == 1992 && local_vf_active == 1) port_count[1992]++; 
              else if (local_pf_num == 0 && local_vf_num == 1993 && local_vf_active == 1) port_count[1993]++; 
              else if (local_pf_num == 0 && local_vf_num == 1994 && local_vf_active == 1) port_count[1994]++; 
              else if (local_pf_num == 0 && local_vf_num == 1995 && local_vf_active == 1) port_count[1995]++; 
              else if (local_pf_num == 0 && local_vf_num == 1996 && local_vf_active == 1) port_count[1996]++; 
              else if (local_pf_num == 0 && local_vf_num == 1997 && local_vf_active == 1) port_count[1997]++; 
              else if (local_pf_num == 0 && local_vf_num == 1998 && local_vf_active == 1) port_count[1998]++; 
              else if (local_pf_num == 0 && local_vf_num == 1999 && local_vf_active == 1) port_count[1999]++; 
              else if (local_pf_num == 0 && local_vf_num == 2000 && local_vf_active == 1) port_count[2000]++; 
              else if (local_pf_num == 0 && local_vf_num == 2001 && local_vf_active == 1) port_count[2001]++; 
              else if (local_pf_num == 0 && local_vf_num == 2002 && local_vf_active == 1) port_count[2002]++; 
              else if (local_pf_num == 0 && local_vf_num == 2003 && local_vf_active == 1) port_count[2003]++; 
              else if (local_pf_num == 0 && local_vf_num == 2004 && local_vf_active == 1) port_count[2004]++; 
              else if (local_pf_num == 0 && local_vf_num == 2005 && local_vf_active == 1) port_count[2005]++; 
              else if (local_pf_num == 0 && local_vf_num == 2006 && local_vf_active == 1) port_count[2006]++; 
              else if (local_pf_num == 0 && local_vf_num == 2007 && local_vf_active == 1) port_count[2007]++; 
              else if (local_pf_num == 0 && local_vf_num == 2008 && local_vf_active == 1) port_count[2008]++; 
              else if (local_pf_num == 0 && local_vf_num == 2009 && local_vf_active == 1) port_count[2009]++; 
              else if (local_pf_num == 0 && local_vf_num == 2010 && local_vf_active == 1) port_count[2010]++; 
              else if (local_pf_num == 0 && local_vf_num == 2011 && local_vf_active == 1) port_count[2011]++; 
              else if (local_pf_num == 0 && local_vf_num == 2012 && local_vf_active == 1) port_count[2012]++; 
              else if (local_pf_num == 0 && local_vf_num == 2013 && local_vf_active == 1) port_count[2013]++; 
              else if (local_pf_num == 0 && local_vf_num == 2014 && local_vf_active == 1) port_count[2014]++; 
              else if (local_pf_num == 0 && local_vf_num == 2015 && local_vf_active == 1) port_count[2015]++; 
              else if (local_pf_num == 0 && local_vf_num == 2016 && local_vf_active == 1) port_count[2016]++; 
              else if (local_pf_num == 0 && local_vf_num == 2017 && local_vf_active == 1) port_count[2017]++; 
              else if (local_pf_num == 0 && local_vf_num == 2018 && local_vf_active == 1) port_count[2018]++; 
              else if (local_pf_num == 0 && local_vf_num == 2019 && local_vf_active == 1) port_count[2019]++; 
              else if (local_pf_num == 0 && local_vf_num == 2020 && local_vf_active == 1) port_count[2020]++; 
              else if (local_pf_num == 0 && local_vf_num == 2021 && local_vf_active == 1) port_count[2021]++; 
              else if (local_pf_num == 0 && local_vf_num == 2022 && local_vf_active == 1) port_count[2022]++; 
              else if (local_pf_num == 0 && local_vf_num == 2023 && local_vf_active == 1) port_count[2023]++; 
              else if (local_pf_num == 0 && local_vf_num == 2024 && local_vf_active == 1) port_count[2024]++; 
              else if (local_pf_num == 0 && local_vf_num == 2025 && local_vf_active == 1) port_count[2025]++; 
              else if (local_pf_num == 0 && local_vf_num == 2026 && local_vf_active == 1) port_count[2026]++; 
              else if (local_pf_num == 0 && local_vf_num == 2027 && local_vf_active == 1) port_count[2027]++; 
              else if (local_pf_num == 0 && local_vf_num == 2028 && local_vf_active == 1) port_count[2028]++; 
              else if (local_pf_num == 0 && local_vf_num == 2029 && local_vf_active == 1) port_count[2029]++; 
              else if (local_pf_num == 0 && local_vf_num == 2030 && local_vf_active == 1) port_count[2030]++; 
              else if (local_pf_num == 0 && local_vf_num == 2031 && local_vf_active == 1) port_count[2031]++; 
              else if (local_pf_num == 0 && local_vf_num == 2032 && local_vf_active == 1) port_count[2032]++; 
              else if (local_pf_num == 0 && local_vf_num == 2033 && local_vf_active == 1) port_count[2033]++; 
              else if (local_pf_num == 0 && local_vf_num == 2034 && local_vf_active == 1) port_count[2034]++; 
              else if (local_pf_num == 0 && local_vf_num == 2035 && local_vf_active == 1) port_count[2035]++; 
              else if (local_pf_num == 0 && local_vf_num == 2036 && local_vf_active == 1) port_count[2036]++; 
              else if (local_pf_num == 0 && local_vf_num == 2037 && local_vf_active == 1) port_count[2037]++; 
              else if (local_pf_num == 0 && local_vf_num == 2038 && local_vf_active == 1) port_count[2038]++; 
              else if (local_pf_num == 0 && local_vf_num == 2039 && local_vf_active == 1) port_count[2039]++; 
              else if (local_pf_num == 0 && local_vf_num == 2040 && local_vf_active == 1) port_count[2040]++; 
              else if (local_pf_num == 0 && local_vf_num == 2041 && local_vf_active == 1) port_count[2041]++; 
              else if (local_pf_num == 0 && local_vf_num == 2042 && local_vf_active == 1) port_count[2042]++; 
              else if (local_pf_num == 0 && local_vf_num == 2043 && local_vf_active == 1) port_count[2043]++; 
              else if (local_pf_num == 0 && local_vf_num == 2044 && local_vf_active == 1) port_count[2044]++; 
              else if (local_pf_num == 0 && local_vf_num == 2045 && local_vf_active == 1) port_count[2045]++; 
              else if (local_pf_num == 0 && local_vf_num == 2046 && local_vf_active == 1) port_count[2046]++; 
              else if (local_pf_num == 0 && local_vf_num == 2047 && local_vf_active == 1) port_count[2047]++; 
              `endif

              for(int j=0; j < (local_tlp_length*32); j++) local_my_payload[j] = 1'b1;
              local_payload = (random_value) & local_my_payload;
              `uvm_info("body", $sformatf("TLP Length = %h and Payload = %h and Random Value generated = %h",local_tlp_length,local_payload,random_value), UVM_LOW)
              //=============================================
              // Starting request sequence on Host master
              //=============================================
              `uvm_do_on_with(master_seq_1, p_sequencer.master_sequencer_H, { tlp_length  == local_tlp_length  ;
                                                                               pf_num      == local_pf_num      ;
                                                                               vf_num      == local_vf_num      ;
                                                                               vf_active   == local_vf_active   ;
                                                                               payload     == local_payload     ;
                                                                               direction   == 1'b0              ;
                                                                            })
               //end
          end
          /////////////////////////////////////////////////////
          //DEVICE TO HOST
          /////////////////////////////////////////////////////
     `ifndef TB_CONFIG_4
          begin
             
            `payload_generate('h0,'h0,'h0);

            `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D0, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                      
                                                                                              })
          end
          begin
             
            `payload_generate('h1,'h0,'h0);

            `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                      
                                                                                              })
          end
         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h2,'h0,'h0);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D2, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h3,'h0,'h0);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D3, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                     
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h4,'h0,'h0);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D4, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                     
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h5,'h0,'h0);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D5, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                     
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h6,'h0,'h0);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D6, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                      
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h7,'h0,'h0);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D7, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                      
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h0,'h0,'h1);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D8, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                    
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h1,'h0,'h1);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D9, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h2,'h0,'h1);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D10, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                     
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h3,'h0,'h1);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D11, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                    
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h4,'h0,'h1);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D12, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                   
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h5,'h0,'h1);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D13, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                      
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h6,'h0,'h1);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D14, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                      
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h7,'h0,'h1);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D15, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                      
                                                                                              })
           

         end
         `ifdef TB_CONFIG_2
         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h0,'h7FF,'h1);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_DN0, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                      
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h1,'h7FF,'h1);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_DN1, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                      
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h2,'h7FF,'h1);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_DN2, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                      
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h3,'h7FF,'h1);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_DN3, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                      
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h4,'h7FF,'h1);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_DN4, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                      
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h5,'h7FF,'h1);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_DN5, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                      
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h6,'h7FF,'h1);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_DN6, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                      
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h7,'h7FF,'h1);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_DN7, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                      
                                                                                              })
           

         end
         `endif

         `ifdef TB_CONFIG_3
        begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h0,'h7FF,'h1);

          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_DN0, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                      
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h1,'h7FF,'h1);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_DN1, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                      
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h2,'h7FF,'h1);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_DN2, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                      
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h3,'h7FF,'h1);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_DN3, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                      
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h4,'h7FF,'h1);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_DN4, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                      
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h5,'h7FF,'h1);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_DN5, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                      
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h6,'h7FF,'h1);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_DN6, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                      
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h7,'h7FF,'h1);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_DN7, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                      
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h0,`RANDOM_VF,'h1);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_DN8, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                      
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h1,`RANDOM_VF,'h1);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_DN9, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                      
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h2,`RANDOM_VF,'h1);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_DN10, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                      
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h3,`RANDOM_VF,'h1);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_DN11, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                      
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h4,`RANDOM_VF,'h1);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_DN12, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                      
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h5,`RANDOM_VF,'h1);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_DN13, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                      
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h6,`RANDOM_VF,'h1);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_DN14, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                      
                                                                                              })
           

         end

         begin
          //===============================================
          // Generating the payload w.r.t TLP length field
          //===============================================

          `payload_generate('h7,`RANDOM_VF,'h1);
 
          //=============================================
          // Starting request sequence on Host master
          //=============================================
          
         
         `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_DN15, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                      
                                                                                              })
           

         end
         `endif
      `endif
       
      `ifdef TB_CONFIG_4
        `payload_generate('h0,0,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D0, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,2,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D2, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,3,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D3, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,4,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D4, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,5,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D5, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,6,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D6, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,7,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D7, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,8,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D8, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,9,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D9, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,10,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D10, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,11,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D11, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,12,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D12, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,13,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D13, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,14,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D14, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,15,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D15, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,16,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D16, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,17,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D17, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,18,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D18, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,19,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D19, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,20,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D20, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,21,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D21, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,22,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D22, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,23,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D23, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,24,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D24, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,25,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D25, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,26,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D26, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,27,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D27, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,28,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D28, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,29,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D29, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,30,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D30, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,31,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D31, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,32,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D32, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,33,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D33, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,34,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D34, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,35,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D35, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,36,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D36, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,37,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D37, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,38,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D38, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,39,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D39, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,40,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D40, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,41,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D41, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,42,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D42, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,43,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D43, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,44,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D44, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,45,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D45, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,46,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D46, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,47,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D47, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,48,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D48, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,49,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D49, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,50,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D50, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,51,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D51, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,52,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D52, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,53,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D53, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,54,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D54, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,55,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D55, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,56,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D56, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,57,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D57, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,58,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D58, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,59,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D59, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,60,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D60, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,61,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D61, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,62,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D62, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,63,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D63, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,64,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D64, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,65,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D65, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,66,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D66, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,67,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D67, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,68,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D68, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,69,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D69, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,70,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D70, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,71,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D71, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,72,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D72, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,73,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D73, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,74,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D74, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,75,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D75, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,76,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D76, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,77,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D77, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,78,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D78, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,79,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D79, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,80,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D80, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,81,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D81, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,82,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D82, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,83,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D83, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,84,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D84, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,85,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D85, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,86,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D86, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,87,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D87, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,88,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D88, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,89,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D89, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,90,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D90, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,91,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D91, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,92,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D92, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,93,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D93, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,94,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D94, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,95,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D95, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,96,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D96, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,97,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D97, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,98,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D98, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,99,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D99, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,100,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D100, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,101,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D101, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,102,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D102, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,103,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D103, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,104,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D104, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,105,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D105, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,106,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D106, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,107,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D107, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,108,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D108, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,109,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D109, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,110,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D110, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,111,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D111, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,112,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D112, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,113,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D113, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,114,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D114, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,115,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D115, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,116,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D116, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,117,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D117, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,118,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D118, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,119,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D119, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,120,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D120, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,121,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D121, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,122,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D122, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,123,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D123, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,124,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D124, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,125,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D125, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,126,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D126, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,127,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D127, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,128,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D128, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,129,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D129, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,130,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D130, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,131,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D131, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,132,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D132, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,133,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D133, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,134,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D134, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,135,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D135, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,136,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D136, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,137,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D137, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,138,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D138, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,139,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D139, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,140,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D140, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,141,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D141, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,142,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D142, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,143,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D143, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,144,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D144, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,145,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D145, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,146,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D146, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,147,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D147, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,148,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D148, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,149,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D149, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,150,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D150, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,151,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D151, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,152,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D152, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,153,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D153, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,154,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D154, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,155,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D155, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,156,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D156, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,157,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D157, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,158,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D158, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,159,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D159, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,160,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D160, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,161,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D161, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,162,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D162, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,163,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D163, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,164,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D164, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,165,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D165, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,166,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D166, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,167,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D167, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,168,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D168, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,169,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D169, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,170,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D170, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,171,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D171, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,172,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D172, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,173,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D173, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,174,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D174, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,175,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D175, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,176,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D176, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,177,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D177, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,178,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D178, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,179,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D179, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,180,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D180, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,181,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D181, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,182,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D182, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,183,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D183, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,184,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D184, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,185,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D185, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,186,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D186, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,187,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D187, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,188,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D188, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,189,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D189, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,190,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D190, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,191,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D191, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,192,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D192, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,193,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D193, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,194,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D194, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,195,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D195, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,196,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D196, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,197,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D197, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,198,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D198, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,199,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D199, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,200,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D200, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,201,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D201, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,202,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D202, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,203,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D203, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,204,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D204, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,205,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D205, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,206,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D206, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,207,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D207, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,208,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D208, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,209,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D209, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,210,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D210, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,211,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D211, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,212,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D212, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,213,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D213, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,214,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D214, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,215,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D215, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,216,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D216, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,217,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D217, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,218,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D218, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,219,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D219, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,220,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D220, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,221,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D221, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,222,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D222, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,223,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D223, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,224,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D224, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,225,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D225, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,226,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D226, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,227,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D227, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,228,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D228, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,229,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D229, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,230,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D230, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,231,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D231, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,232,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D232, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,233,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D233, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,234,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D234, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,235,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D235, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,236,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D236, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,237,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D237, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,238,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D238, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,239,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D239, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,240,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D240, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,241,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D241, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,242,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D242, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,243,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D243, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,244,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D244, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,245,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D245, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,246,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D246, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,247,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D247, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,248,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D248, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,249,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D249, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,250,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D250, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,251,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D251, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,252,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D252, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,253,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D253, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,254,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D254, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,255,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D255, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,256,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D256, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,257,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D257, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,258,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D258, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,259,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D259, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,260,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D260, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,261,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D261, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,262,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D262, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,263,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D263, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,264,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D264, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,265,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D265, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,266,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D266, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,267,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D267, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,268,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D268, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,269,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D269, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,270,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D270, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,271,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D271, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,272,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D272, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,273,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D273, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,274,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D274, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,275,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D275, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,276,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D276, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,277,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D277, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,278,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D278, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,279,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D279, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,280,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D280, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,281,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D281, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,282,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D282, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,283,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D283, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,284,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D284, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,285,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D285, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,286,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D286, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,287,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D287, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,288,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D288, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,289,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D289, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,290,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D290, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,291,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D291, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,292,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D292, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,293,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D293, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,294,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D294, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,295,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D295, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,296,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D296, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,297,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D297, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,298,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D298, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,299,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D299, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,300,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D300, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,301,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D301, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,302,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D302, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,303,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D303, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,304,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D304, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,305,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D305, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,306,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D306, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,307,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D307, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,308,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D308, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,309,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D309, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,310,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D310, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,311,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D311, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,312,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D312, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,313,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D313, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,314,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D314, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,315,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D315, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,316,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D316, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,317,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D317, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,318,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D318, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,319,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D319, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,320,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D320, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,321,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D321, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,322,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D322, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,323,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D323, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,324,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D324, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,325,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D325, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,326,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D326, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,327,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D327, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,328,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D328, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,329,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D329, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,330,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D330, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,331,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D331, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,332,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D332, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,333,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D333, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,334,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D334, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,335,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D335, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,336,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D336, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,337,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D337, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,338,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D338, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,339,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D339, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,340,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D340, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,341,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D341, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,342,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D342, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,343,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D343, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,344,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D344, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,345,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D345, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,346,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D346, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,347,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D347, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,348,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D348, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,349,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D349, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,350,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D350, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,351,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D351, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,352,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D352, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,353,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D353, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,354,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D354, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,355,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D355, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,356,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D356, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,357,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D357, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,358,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D358, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,359,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D359, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,360,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D360, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,361,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D361, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,362,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D362, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,363,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D363, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,364,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D364, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,365,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D365, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,366,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D366, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,367,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D367, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,368,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D368, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,369,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D369, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,370,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D370, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,371,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D371, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,372,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D372, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,373,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D373, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,374,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D374, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,375,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D375, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,376,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D376, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,377,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D377, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,378,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D378, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,379,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D379, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,380,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D380, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,381,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D381, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,382,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D382, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,383,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D383, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,384,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D384, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,385,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D385, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,386,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D386, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,387,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D387, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,388,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D388, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,389,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D389, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,390,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D390, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,391,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D391, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,392,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D392, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,393,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D393, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,394,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D394, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,395,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D395, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,396,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D396, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,397,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D397, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,398,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D398, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,399,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D399, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,400,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D400, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,401,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D401, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,402,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D402, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,403,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D403, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,404,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D404, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,405,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D405, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,406,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D406, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,407,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D407, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,408,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D408, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,409,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D409, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,410,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D410, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,411,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D411, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,412,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D412, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,413,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D413, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,414,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D414, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,415,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D415, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,416,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D416, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,417,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D417, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,418,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D418, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,419,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D419, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,420,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D420, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,421,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D421, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,422,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D422, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,423,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D423, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,424,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D424, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,425,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D425, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,426,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D426, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,427,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D427, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,428,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D428, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,429,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D429, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,430,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D430, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,431,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D431, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,432,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D432, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,433,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D433, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,434,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D434, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,435,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D435, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,436,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D436, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,437,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D437, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,438,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D438, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,439,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D439, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,440,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D440, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,441,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D441, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,442,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D442, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,443,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D443, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,444,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D444, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,445,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D445, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,446,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D446, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,447,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D447, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,448,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D448, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,449,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D449, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,450,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D450, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,451,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D451, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,452,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D452, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,453,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D453, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,454,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D454, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,455,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D455, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,456,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D456, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,457,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D457, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,458,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D458, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,459,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D459, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,460,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D460, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,461,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D461, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,462,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D462, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,463,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D463, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,464,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D464, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,465,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D465, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,466,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D466, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,467,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D467, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,468,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D468, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,469,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D469, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,470,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D470, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,471,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D471, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,472,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D472, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,473,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D473, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,474,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D474, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,475,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D475, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,476,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D476, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,477,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D477, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,478,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D478, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,479,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D479, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,480,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D480, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,481,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D481, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,482,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D482, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,483,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D483, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,484,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D484, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,485,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D485, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,486,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D486, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,487,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D487, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,488,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D488, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,489,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D489, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,490,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D490, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,491,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D491, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,492,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D492, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,493,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D493, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,494,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D494, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,495,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D495, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,496,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D496, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,497,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D497, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,498,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D498, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,499,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D499, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,500,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D500, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,501,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D501, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,502,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D502, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,503,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D503, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,504,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D504, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,505,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D505, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,506,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D506, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,507,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D507, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,508,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D508, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,509,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D509, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,510,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D510, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,511,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D511, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,512,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D512, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,513,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D513, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,514,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D514, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,515,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D515, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,516,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D516, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,517,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D517, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,518,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D518, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,519,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D519, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,520,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D520, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,521,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D521, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,522,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D522, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,523,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D523, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,524,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D524, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,525,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D525, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,526,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D526, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,527,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D527, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,528,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D528, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,529,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D529, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,530,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D530, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,531,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D531, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,532,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D532, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,533,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D533, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,534,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D534, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,535,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D535, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,536,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D536, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,537,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D537, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,538,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D538, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,539,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D539, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,540,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D540, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,541,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D541, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,542,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D542, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,543,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D543, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,544,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D544, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,545,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D545, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,546,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D546, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,547,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D547, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,548,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D548, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,549,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D549, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,550,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D550, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,551,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D551, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,552,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D552, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,553,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D553, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,554,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D554, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,555,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D555, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,556,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D556, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,557,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D557, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,558,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D558, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,559,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D559, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,560,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D560, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,561,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D561, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,562,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D562, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,563,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D563, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,564,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D564, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,565,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D565, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,566,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D566, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,567,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D567, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,568,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D568, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,569,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D569, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,570,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D570, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,571,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D571, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,572,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D572, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,573,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D573, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,574,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D574, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,575,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D575, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,576,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D576, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,577,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D577, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,578,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D578, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,579,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D579, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,580,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D580, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,581,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D581, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,582,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D582, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,583,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D583, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,584,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D584, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,585,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D585, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,586,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D586, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,587,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D587, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,588,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D588, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,589,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D589, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,590,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D590, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,591,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D591, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,592,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D592, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,593,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D593, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,594,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D594, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,595,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D595, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,596,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D596, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,597,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D597, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,598,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D598, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,599,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D599, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,600,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D600, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,601,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D601, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,602,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D602, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,603,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D603, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,604,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D604, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,605,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D605, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,606,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D606, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,607,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D607, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,608,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D608, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,609,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D609, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,610,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D610, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,611,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D611, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,612,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D612, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,613,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D613, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,614,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D614, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,615,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D615, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,616,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D616, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,617,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D617, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,618,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D618, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,619,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D619, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,620,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D620, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,621,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D621, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,622,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D622, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,623,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D623, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,624,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D624, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,625,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D625, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,626,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D626, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,627,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D627, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,628,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D628, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,629,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D629, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,630,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D630, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,631,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D631, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,632,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D632, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,633,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D633, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,634,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D634, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,635,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D635, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,636,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D636, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,637,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D637, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,638,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D638, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,639,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D639, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,640,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D640, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,641,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D641, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,642,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D642, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,643,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D643, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,644,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D644, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,645,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D645, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,646,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D646, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,647,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D647, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,648,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D648, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,649,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D649, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,650,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D650, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,651,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D651, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,652,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D652, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,653,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D653, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,654,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D654, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,655,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D655, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,656,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D656, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,657,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D657, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,658,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D658, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,659,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D659, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,660,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D660, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,661,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D661, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,662,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D662, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,663,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D663, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,664,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D664, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,665,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D665, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,666,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D666, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,667,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D667, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,668,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D668, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,669,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D669, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,670,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D670, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,671,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D671, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,672,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D672, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,673,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D673, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,674,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D674, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,675,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D675, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,676,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D676, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,677,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D677, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,678,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D678, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,679,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D679, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,680,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D680, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,681,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D681, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,682,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D682, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,683,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D683, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,684,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D684, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,685,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D685, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,686,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D686, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,687,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D687, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,688,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D688, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,689,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D689, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,690,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D690, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,691,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D691, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,692,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D692, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,693,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D693, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,694,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D694, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,695,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D695, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,696,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D696, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,697,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D697, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,698,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D698, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,699,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D699, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,700,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D700, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,701,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D701, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,702,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D702, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,703,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D703, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,704,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D704, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,705,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D705, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,706,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D706, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,707,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D707, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,708,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D708, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,709,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D709, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,710,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D710, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,711,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D711, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,712,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D712, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,713,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D713, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,714,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D714, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,715,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D715, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,716,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D716, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,717,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D717, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,718,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D718, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,719,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D719, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,720,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D720, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,721,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D721, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,722,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D722, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,723,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D723, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,724,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D724, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,725,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D725, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,726,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D726, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,727,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D727, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,728,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D728, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,729,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D729, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,730,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D730, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,731,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D731, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,732,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D732, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,733,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D733, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,734,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D734, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,735,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D735, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,736,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D736, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,737,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D737, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,738,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D738, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,739,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D739, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,740,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D740, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,741,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D741, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,742,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D742, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,743,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D743, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,744,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D744, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,745,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D745, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,746,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D746, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,747,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D747, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,748,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D748, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,749,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D749, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,750,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D750, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,751,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D751, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,752,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D752, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,753,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D753, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,754,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D754, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,755,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D755, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,756,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D756, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,757,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D757, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,758,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D758, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,759,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D759, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,760,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D760, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,761,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D761, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,762,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D762, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,763,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D763, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,764,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D764, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,765,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D765, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,766,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D766, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,767,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D767, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,768,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D768, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,769,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D769, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,770,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D770, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,771,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D771, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,772,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D772, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,773,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D773, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,774,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D774, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,775,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D775, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,776,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D776, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,777,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D777, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,778,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D778, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,779,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D779, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,780,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D780, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,781,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D781, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,782,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D782, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,783,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D783, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,784,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D784, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,785,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D785, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,786,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D786, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,787,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D787, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,788,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D788, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,789,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D789, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,790,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D790, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,791,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D791, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,792,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D792, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,793,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D793, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,794,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D794, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,795,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D795, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,796,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D796, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,797,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D797, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,798,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D798, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,799,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D799, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,800,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D800, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,801,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D801, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,802,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D802, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,803,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D803, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,804,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D804, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,805,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D805, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,806,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D806, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,807,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D807, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,808,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D808, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,809,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D809, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,810,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D810, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,811,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D811, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,812,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D812, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,813,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D813, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,814,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D814, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,815,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D815, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,816,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D816, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,817,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D817, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,818,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D818, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,819,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D819, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,820,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D820, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,821,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D821, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,822,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D822, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,823,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D823, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,824,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D824, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,825,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D825, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,826,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D826, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,827,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D827, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,828,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D828, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,829,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D829, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,830,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D830, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,831,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D831, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,832,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D832, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,833,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D833, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,834,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D834, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,835,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D835, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,836,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D836, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,837,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D837, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,838,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D838, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,839,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D839, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,840,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D840, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,841,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D841, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,842,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D842, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,843,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D843, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,844,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D844, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,845,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D845, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,846,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D846, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,847,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D847, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,848,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D848, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,849,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D849, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,850,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D850, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,851,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D851, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,852,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D852, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,853,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D853, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,854,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D854, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,855,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D855, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,856,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D856, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,857,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D857, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,858,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D858, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,859,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D859, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,860,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D860, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,861,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D861, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,862,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D862, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,863,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D863, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,864,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D864, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,865,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D865, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,866,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D866, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,867,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D867, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,868,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D868, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,869,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D869, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,870,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D870, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,871,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D871, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,872,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D872, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,873,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D873, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,874,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D874, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,875,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D875, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,876,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D876, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,877,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D877, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,878,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D878, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,879,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D879, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,880,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D880, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,881,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D881, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,882,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D882, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,883,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D883, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,884,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D884, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,885,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D885, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,886,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D886, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,887,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D887, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,888,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D888, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,889,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D889, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,890,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D890, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,891,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D891, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,892,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D892, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,893,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D893, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,894,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D894, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,895,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D895, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,896,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D896, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,897,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D897, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,898,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D898, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,899,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D899, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,900,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D900, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,901,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D901, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,902,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D902, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,903,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D903, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,904,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D904, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,905,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D905, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,906,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D906, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,907,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D907, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,908,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D908, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,909,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D909, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,910,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D910, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,911,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D911, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,912,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D912, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,913,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D913, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,914,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D914, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,915,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D915, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,916,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D916, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,917,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D917, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,918,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D918, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,919,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D919, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,920,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D920, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,921,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D921, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,922,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D922, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,923,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D923, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,924,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D924, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,925,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D925, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,926,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D926, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,927,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D927, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,928,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D928, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,929,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D929, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,930,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D930, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,931,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D931, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,932,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D932, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,933,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D933, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,934,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D934, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,935,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D935, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,936,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D936, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,937,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D937, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,938,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D938, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,939,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D939, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,940,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D940, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,941,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D941, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,942,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D942, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,943,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D943, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,944,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D944, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,945,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D945, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,946,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D946, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,947,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D947, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,948,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D948, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,949,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D949, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,950,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D950, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,951,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D951, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,952,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D952, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,953,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D953, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,954,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D954, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,955,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D955, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,956,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D956, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,957,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D957, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,958,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D958, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,959,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D959, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,960,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D960, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,961,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D961, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,962,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D962, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,963,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D963, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,964,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D964, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,965,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D965, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,966,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D966, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,967,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D967, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,968,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D968, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,969,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D969, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,970,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D970, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,971,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D971, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,972,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D972, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,973,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D973, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,974,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D974, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,975,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D975, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,976,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D976, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,977,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D977, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,978,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D978, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,979,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D979, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,980,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D980, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,981,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D981, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,982,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D982, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,983,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D983, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,984,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D984, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,985,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D985, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,986,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D986, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,987,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D987, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,988,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D988, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,989,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D989, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,990,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D990, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,991,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D991, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,992,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D992, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,993,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D993, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,994,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D994, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,995,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D995, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,996,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D996, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,997,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D997, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,998,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D998, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,999,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D999, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1000,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1000, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1001,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1001, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1002,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1002, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1003,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1003, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1004,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1004, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1005,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1005, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1006,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1006, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1007,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1007, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1008,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1008, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1009,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1009, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1010,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1010, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1011,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1011, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1012,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1012, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1013,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1013, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1014,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1014, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1015,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1015, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1016,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1016, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1017,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1017, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1018,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1018, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1019,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1019, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1020,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1020, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1021,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1021, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1022,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1022, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1023,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1023, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1024,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1024, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1025,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1025, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1026,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1026, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1027,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1027, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1028,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1028, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1029,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1029, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1030,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1030, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1031,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1031, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1032,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1032, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1033,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1033, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1034,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1034, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1035,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1035, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1036,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1036, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1037,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1037, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1038,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1038, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1039,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1039, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1040,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1040, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1041,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1041, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1042,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1042, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1043,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1043, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1044,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1044, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1045,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1045, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1046,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1046, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1047,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1047, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1048,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1048, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1049,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1049, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1050,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1050, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1051,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1051, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1052,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1052, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1053,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1053, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1054,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1054, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1055,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1055, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1056,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1056, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1057,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1057, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1058,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1058, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1059,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1059, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1060,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1060, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1061,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1061, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1062,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1062, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1063,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1063, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1064,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1064, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1065,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1065, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1066,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1066, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1067,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1067, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1068,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1068, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1069,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1069, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1070,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1070, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1071,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1071, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1072,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1072, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1073,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1073, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1074,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1074, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1075,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1075, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1076,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1076, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1077,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1077, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1078,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1078, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1079,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1079, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1080,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1080, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1081,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1081, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1082,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1082, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1083,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1083, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1084,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1084, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1085,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1085, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1086,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1086, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1087,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1087, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1088,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1088, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1089,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1089, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1090,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1090, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1091,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1091, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1092,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1092, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1093,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1093, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1094,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1094, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1095,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1095, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1096,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1096, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1097,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1097, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1098,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1098, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1099,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1099, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1100,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1100, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1101,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1101, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1102,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1102, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1103,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1103, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1104,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1104, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1105,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1105, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1106,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1106, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1107,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1107, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1108,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1108, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1109,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1109, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1110,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1110, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1111,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1111, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1112,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1112, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1113,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1113, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1114,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1114, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1115,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1115, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1116,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1116, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1117,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1117, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1118,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1118, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1119,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1119, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1120,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1120, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1121,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1121, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1122,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1122, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1123,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1123, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1124,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1124, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1125,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1125, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1126,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1126, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1127,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1127, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1128,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1128, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1129,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1129, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1130,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1130, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1131,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1131, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1132,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1132, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1133,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1133, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1134,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1134, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1135,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1135, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1136,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1136, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1137,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1137, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1138,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1138, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1139,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1139, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1140,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1140, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1141,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1141, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1142,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1142, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1143,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1143, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1144,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1144, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1145,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1145, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1146,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1146, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1147,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1147, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1148,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1148, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1149,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1149, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1150,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1150, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1151,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1151, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1152,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1152, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1153,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1153, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1154,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1154, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1155,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1155, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1156,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1156, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1157,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1157, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1158,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1158, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1159,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1159, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1160,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1160, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1161,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1161, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1162,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1162, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1163,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1163, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1164,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1164, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1165,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1165, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1166,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1166, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1167,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1167, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1168,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1168, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1169,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1169, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1170,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1170, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1171,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1171, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1172,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1172, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1173,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1173, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1174,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1174, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1175,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1175, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1176,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1176, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1177,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1177, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1178,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1178, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1179,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1179, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1180,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1180, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1181,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1181, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1182,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1182, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1183,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1183, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1184,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1184, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1185,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1185, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1186,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1186, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1187,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1187, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1188,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1188, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1189,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1189, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1190,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1190, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1191,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1191, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1192,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1192, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1193,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1193, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1194,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1194, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1195,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1195, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1196,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1196, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1197,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1197, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1198,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1198, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1199,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1199, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1200,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1200, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1201,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1201, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1202,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1202, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1203,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1203, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1204,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1204, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1205,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1205, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1206,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1206, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1207,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1207, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1208,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1208, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1209,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1209, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1210,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1210, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1211,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1211, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1212,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1212, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1213,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1213, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1214,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1214, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1215,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1215, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1216,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1216, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1217,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1217, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1218,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1218, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1219,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1219, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1220,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1220, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1221,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1221, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1222,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1222, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1223,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1223, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1224,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1224, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1225,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1225, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1226,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1226, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1227,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1227, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1228,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1228, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1229,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1229, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1230,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1230, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1231,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1231, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1232,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1232, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1233,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1233, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1234,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1234, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1235,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1235, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1236,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1236, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1237,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1237, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1238,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1238, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1239,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1239, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1240,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1240, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1241,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1241, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1242,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1242, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1243,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1243, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1244,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1244, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1245,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1245, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1246,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1246, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1247,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1247, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1248,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1248, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1249,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1249, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1250,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1250, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1251,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1251, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1252,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1252, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1253,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1253, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1254,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1254, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1255,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1255, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1256,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1256, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1257,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1257, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1258,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1258, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1259,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1259, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1260,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1260, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1261,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1261, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1262,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1262, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1263,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1263, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1264,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1264, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1265,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1265, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1266,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1266, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1267,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1267, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1268,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1268, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1269,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1269, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1270,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1270, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1271,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1271, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1272,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1272, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1273,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1273, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1274,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1274, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1275,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1275, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1276,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1276, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1277,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1277, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1278,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1278, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1279,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1279, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1280,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1280, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1281,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1281, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1282,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1282, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1283,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1283, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1284,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1284, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1285,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1285, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1286,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1286, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1287,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1287, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1288,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1288, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1289,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1289, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1290,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1290, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1291,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1291, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1292,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1292, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1293,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1293, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1294,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1294, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1295,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1295, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1296,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1296, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1297,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1297, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1298,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1298, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1299,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1299, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1300,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1300, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1301,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1301, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1302,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1302, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1303,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1303, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1304,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1304, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1305,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1305, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1306,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1306, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1307,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1307, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1308,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1308, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1309,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1309, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1310,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1310, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1311,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1311, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1312,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1312, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1313,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1313, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1314,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1314, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1315,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1315, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1316,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1316, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1317,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1317, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1318,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1318, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1319,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1319, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1320,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1320, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1321,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1321, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1322,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1322, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1323,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1323, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1324,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1324, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1325,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1325, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1326,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1326, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1327,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1327, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1328,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1328, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1329,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1329, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1330,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1330, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1331,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1331, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1332,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1332, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1333,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1333, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1334,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1334, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1335,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1335, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1336,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1336, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1337,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1337, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1338,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1338, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1339,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1339, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1340,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1340, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1341,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1341, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1342,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1342, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1343,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1343, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1344,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1344, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1345,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1345, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1346,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1346, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1347,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1347, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1348,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1348, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1349,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1349, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1350,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1350, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1351,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1351, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1352,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1352, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1353,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1353, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1354,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1354, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1355,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1355, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1356,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1356, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1357,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1357, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1358,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1358, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1359,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1359, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1360,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1360, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1361,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1361, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1362,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1362, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1363,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1363, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1364,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1364, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1365,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1365, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1366,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1366, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1367,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1367, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1368,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1368, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1369,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1369, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1370,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1370, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1371,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1371, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1372,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1372, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1373,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1373, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1374,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1374, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1375,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1375, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1376,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1376, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1377,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1377, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1378,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1378, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1379,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1379, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1380,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1380, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1381,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1381, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1382,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1382, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1383,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1383, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1384,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1384, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1385,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1385, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1386,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1386, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1387,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1387, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1388,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1388, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1389,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1389, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1390,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1390, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1391,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1391, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1392,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1392, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1393,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1393, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1394,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1394, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1395,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1395, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1396,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1396, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1397,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1397, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1398,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1398, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1399,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1399, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1400,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1400, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1401,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1401, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1402,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1402, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1403,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1403, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1404,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1404, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1405,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1405, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1406,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1406, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1407,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1407, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1408,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1408, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1409,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1409, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1410,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1410, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1411,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1411, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1412,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1412, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1413,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1413, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1414,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1414, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1415,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1415, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1416,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1416, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1417,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1417, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1418,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1418, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1419,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1419, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1420,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1420, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1421,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1421, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1422,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1422, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1423,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1423, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1424,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1424, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1425,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1425, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1426,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1426, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1427,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1427, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1428,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1428, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1429,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1429, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1430,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1430, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1431,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1431, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1432,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1432, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1433,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1433, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1434,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1434, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1435,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1435, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1436,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1436, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1437,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1437, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1438,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1438, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1439,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1439, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1440,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1440, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1441,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1441, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1442,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1442, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1443,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1443, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1444,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1444, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1445,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1445, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1446,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1446, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1447,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1447, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1448,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1448, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1449,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1449, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1450,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1450, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1451,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1451, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1452,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1452, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1453,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1453, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1454,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1454, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1455,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1455, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1456,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1456, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1457,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1457, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1458,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1458, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1459,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1459, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1460,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1460, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1461,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1461, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1462,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1462, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1463,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1463, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1464,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1464, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1465,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1465, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1466,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1466, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1467,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1467, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1468,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1468, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1469,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1469, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1470,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1470, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1471,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1471, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1472,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1472, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1473,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1473, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1474,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1474, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1475,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1475, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1476,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1476, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1477,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1477, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1478,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1478, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1479,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1479, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1480,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1480, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1481,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1481, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1482,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1482, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1483,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1483, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1484,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1484, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1485,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1485, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1486,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1486, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1487,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1487, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1488,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1488, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1489,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1489, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1490,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1490, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1491,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1491, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1492,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1492, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1493,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1493, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1494,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1494, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1495,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1495, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1496,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1496, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1497,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1497, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1498,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1498, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1499,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1499, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1500,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1500, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1501,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1501, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1502,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1502, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1503,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1503, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1504,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1504, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1505,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1505, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1506,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1506, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1507,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1507, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1508,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1508, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1509,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1509, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1510,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1510, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1511,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1511, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1512,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1512, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1513,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1513, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1514,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1514, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1515,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1515, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1516,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1516, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1517,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1517, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1518,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1518, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1519,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1519, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1520,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1520, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1521,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1521, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1522,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1522, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1523,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1523, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1524,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1524, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1525,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1525, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1526,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1526, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1527,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1527, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1528,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1528, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1529,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1529, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1530,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1530, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1531,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1531, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1532,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1532, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1533,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1533, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1534,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1534, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1535,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1535, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1536,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1536, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1537,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1537, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1538,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1538, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1539,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1539, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1540,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1540, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1541,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1541, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1542,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1542, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1543,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1543, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1544,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1544, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1545,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1545, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1546,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1546, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1547,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1547, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1548,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1548, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1549,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1549, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1550,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1550, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1551,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1551, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1552,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1552, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1553,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1553, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1554,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1554, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1555,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1555, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1556,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1556, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1557,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1557, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1558,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1558, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1559,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1559, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1560,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1560, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1561,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1561, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1562,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1562, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1563,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1563, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1564,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1564, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1565,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1565, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1566,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1566, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1567,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1567, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1568,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1568, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1569,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1569, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1570,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1570, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1571,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1571, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1572,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1572, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1573,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1573, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1574,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1574, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1575,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1575, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1576,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1576, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1577,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1577, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1578,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1578, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1579,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1579, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1580,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1580, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1581,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1581, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1582,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1582, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1583,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1583, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1584,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1584, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1585,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1585, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1586,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1586, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1587,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1587, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1588,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1588, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1589,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1589, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1590,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1590, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1591,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1591, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1592,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1592, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1593,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1593, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1594,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1594, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1595,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1595, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1596,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1596, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1597,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1597, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1598,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1598, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1599,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1599, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1600,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1600, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1601,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1601, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1602,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1602, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1603,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1603, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1604,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1604, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1605,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1605, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1606,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1606, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1607,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1607, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1608,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1608, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1609,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1609, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1610,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1610, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1611,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1611, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1612,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1612, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1613,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1613, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1614,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1614, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1615,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1615, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1616,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1616, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1617,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1617, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1618,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1618, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1619,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1619, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1620,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1620, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1621,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1621, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1622,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1622, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1623,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1623, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1624,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1624, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1625,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1625, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1626,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1626, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1627,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1627, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1628,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1628, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1629,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1629, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1630,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1630, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1631,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1631, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1632,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1632, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1633,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1633, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1634,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1634, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1635,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1635, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1636,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1636, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1637,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1637, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1638,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1638, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1639,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1639, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1640,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1640, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1641,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1641, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1642,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1642, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1643,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1643, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1644,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1644, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1645,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1645, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1646,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1646, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1647,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1647, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1648,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1648, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1649,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1649, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1650,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1650, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1651,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1651, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1652,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1652, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1653,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1653, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1654,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1654, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1655,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1655, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1656,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1656, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1657,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1657, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1658,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1658, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1659,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1659, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1660,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1660, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1661,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1661, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1662,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1662, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1663,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1663, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1664,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1664, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1665,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1665, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1666,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1666, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1667,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1667, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1668,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1668, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1669,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1669, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1670,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1670, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1671,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1671, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1672,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1672, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1673,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1673, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1674,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1674, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1675,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1675, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1676,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1676, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1677,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1677, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1678,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1678, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1679,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1679, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1680,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1680, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1681,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1681, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1682,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1682, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1683,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1683, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1684,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1684, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1685,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1685, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1686,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1686, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1687,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1687, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1688,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1688, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1689,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1689, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1690,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1690, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1691,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1691, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1692,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1692, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1693,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1693, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1694,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1694, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1695,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1695, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1696,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1696, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1697,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1697, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1698,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1698, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1699,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1699, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1700,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1700, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1701,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1701, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1702,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1702, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1703,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1703, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1704,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1704, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1705,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1705, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1706,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1706, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1707,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1707, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1708,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1708, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1709,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1709, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1710,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1710, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1711,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1711, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1712,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1712, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1713,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1713, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1714,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1714, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1715,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1715, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1716,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1716, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1717,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1717, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1718,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1718, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1719,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1719, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1720,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1720, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1721,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1721, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1722,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1722, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1723,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1723, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1724,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1724, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1725,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1725, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1726,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1726, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1727,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1727, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1728,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1728, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1729,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1729, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1730,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1730, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1731,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1731, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1732,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1732, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1733,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1733, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1734,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1734, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1735,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1735, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1736,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1736, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1737,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1737, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1738,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1738, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1739,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1739, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1740,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1740, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1741,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1741, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1742,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1742, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1743,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1743, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1744,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1744, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1745,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1745, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1746,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1746, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1747,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1747, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1748,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1748, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1749,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1749, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1750,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1750, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1751,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1751, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1752,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1752, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1753,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1753, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1754,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1754, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1755,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1755, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1756,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1756, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1757,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1757, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1758,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1758, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1759,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1759, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1760,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1760, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1761,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1761, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1762,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1762, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1763,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1763, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1764,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1764, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1765,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1765, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1766,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1766, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1767,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1767, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1768,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1768, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1769,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1769, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1770,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1770, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1771,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1771, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1772,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1772, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1773,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1773, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1774,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1774, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1775,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1775, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1776,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1776, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1777,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1777, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1778,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1778, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1779,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1779, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1780,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1780, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1781,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1781, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1782,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1782, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1783,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1783, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1784,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1784, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1785,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1785, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1786,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1786, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1787,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1787, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1788,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1788, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1789,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1789, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1790,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1790, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1791,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1791, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1792,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1792, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1793,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1793, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1794,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1794, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1795,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1795, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1796,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1796, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1797,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1797, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1798,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1798, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1799,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1799, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1800,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1800, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1801,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1801, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1802,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1802, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1803,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1803, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1804,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1804, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1805,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1805, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1806,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1806, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1807,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1807, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1808,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1808, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1809,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1809, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1810,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1810, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1811,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1811, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1812,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1812, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1813,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1813, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1814,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1814, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1815,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1815, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1816,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1816, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1817,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1817, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1818,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1818, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1819,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1819, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1820,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1820, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1821,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1821, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1822,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1822, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1823,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1823, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1824,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1824, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1825,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1825, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1826,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1826, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1827,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1827, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1828,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1828, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1829,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1829, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1830,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1830, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1831,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1831, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1832,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1832, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1833,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1833, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1834,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1834, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1835,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1835, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1836,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1836, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1837,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1837, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1838,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1838, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1839,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1839, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1840,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1840, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1841,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1841, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1842,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1842, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1843,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1843, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1844,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1844, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1845,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1845, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1846,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1846, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1847,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1847, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1848,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1848, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1849,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1849, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1850,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1850, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1851,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1851, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1852,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1852, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1853,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1853, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1854,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1854, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1855,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1855, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1856,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1856, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1857,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1857, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1858,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1858, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1859,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1859, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1860,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1860, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1861,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1861, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1862,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1862, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1863,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1863, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1864,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1864, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1865,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1865, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1866,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1866, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1867,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1867, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1868,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1868, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1869,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1869, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1870,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1870, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1871,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1871, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1872,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1872, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1873,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1873, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1874,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1874, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1875,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1875, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1876,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1876, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1877,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1877, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1878,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1878, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1879,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1879, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1880,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1880, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1881,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1881, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1882,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1882, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1883,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1883, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1884,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1884, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1885,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1885, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1886,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1886, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1887,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1887, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1888,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1888, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1889,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1889, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1890,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1890, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1891,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1891, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1892,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1892, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1893,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1893, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1894,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1894, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1895,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1895, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1896,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1896, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1897,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1897, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1898,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1898, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1899,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1899, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1900,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1900, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1901,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1901, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1902,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1902, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1903,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1903, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1904,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1904, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1905,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1905, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1906,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1906, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1907,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1907, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1908,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1908, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1909,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1909, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1910,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1910, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1911,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1911, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1912,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1912, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1913,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1913, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1914,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1914, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1915,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1915, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1916,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1916, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1917,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1917, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1918,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1918, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1919,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1919, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1920,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1920, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1921,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1921, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1922,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1922, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1923,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1923, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1924,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1924, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1925,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1925, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1926,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1926, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1927,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1927, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1928,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1928, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1929,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1929, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1930,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1930, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1931,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1931, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1932,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1932, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1933,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1933, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1934,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1934, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1935,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1935, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1936,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1936, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1937,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1937, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1938,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1938, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1939,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1939, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1940,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1940, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1941,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1941, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1942,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1942, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1943,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1943, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1944,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1944, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1945,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1945, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1946,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1946, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1947,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1947, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1948,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1948, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1949,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1949, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1950,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1950, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1951,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1951, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1952,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1952, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1953,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1953, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1954,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1954, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1955,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1955, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1956,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1956, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1957,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1957, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1958,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1958, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1959,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1959, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1960,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1960, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1961,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1961, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1962,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1962, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1963,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1963, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1964,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1964, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1965,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1965, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1966,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1966, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1967,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1967, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1968,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1968, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1969,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1969, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1970,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1970, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1971,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1971, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1972,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1972, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1973,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1973, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1974,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1974, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1975,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1975, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1976,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1976, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1977,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1977, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1978,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1978, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1979,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1979, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1980,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1980, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1981,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1981, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1982,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1982, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1983,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1983, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1984,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1984, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1985,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1985, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1986,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1986, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1987,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1987, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1988,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1988, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1989,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1989, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1990,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1990, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1991,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1991, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1992,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1992, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1993,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1993, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1994,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1994, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1995,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1995, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1996,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1996, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1997,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1997, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1998,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1998, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,1999,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D1999, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,2000,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D2000, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,2001,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D2001, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,2002,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D2002, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,2003,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D2003, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,2004,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D2004, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,2005,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D2005, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,2006,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D2006, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,2007,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D2007, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,2008,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D2008, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,2009,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D2009, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,2010,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D2010, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,2011,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D2011, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,2012,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D2012, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,2013,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D2013, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,2014,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D2014, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,2015,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D2015, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,2016,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D2016, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,2017,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D2017, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,2018,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D2018, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,2019,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D2019, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,2020,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D2020, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,2021,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D2021, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,2022,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D2022, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,2023,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D2023, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,2024,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D2024, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,2025,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D2025, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,2026,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D2026, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,2027,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D2027, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,2028,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D2028, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,2029,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D2029, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,2030,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D2030, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,2031,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D2031, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,2032,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D2032, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,2033,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D2033, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,2034,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D2034, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,2035,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D2035, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,2036,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D2036, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,2037,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D2037, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,2038,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D2038, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,2039,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D2039, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,2040,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D2040, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,2041,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D2041, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,2042,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D2042, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,2043,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D2043, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,2044,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D2044, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,2045,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D2045, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,2046,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D2046, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
        `payload_generate('h0,2047,'h1);
        `uvm_do_on_with(master_seq_2, p_sequencer.master_sequencer_D2047, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;                                                                                                               })
      `endif

       join
       end    

	     uvm_config_db #(int)::set(null,"*","PORT_0_COUNT",port_count[0]);
	     uvm_config_db #(int)::set(null,"*","PORT_1_COUNT",port_count[1]);
	     uvm_config_db #(int)::set(null,"*","PORT_2_COUNT",port_count[2]);
	     uvm_config_db #(int)::set(null,"*","PORT_3_COUNT",port_count[3]);
	     uvm_config_db #(int)::set(null,"*","PORT_4_COUNT",port_count[4]);
	     uvm_config_db #(int)::set(null,"*","PORT_5_COUNT",port_count[5]);
	     uvm_config_db #(int)::set(null,"*","PORT_6_COUNT",port_count[6]);
	     uvm_config_db #(int)::set(null,"*","PORT_7_COUNT",port_count[7]);
	     uvm_config_db #(int)::set(null,"*","PORT_8_COUNT",port_count[8]);
	     uvm_config_db #(int)::set(null,"*","PORT_9_COUNT",port_count[9]);
	     uvm_config_db #(int)::set(null,"*","PORT_10_COUNT",port_count[10]);
	     uvm_config_db #(int)::set(null,"*","PORT_11_COUNT",port_count[11]);
	     uvm_config_db #(int)::set(null,"*","PORT_12_COUNT",port_count[12]);
	     uvm_config_db #(int)::set(null,"*","PORT_13_COUNT",port_count[13]);
	     uvm_config_db #(int)::set(null,"*","PORT_14_COUNT",port_count[14]);
	     uvm_config_db #(int)::set(null,"*","PORT_15_COUNT",port_count[15]);
	     `ifndef TB_CONFIG_1
       uvm_config_db #(int)::set(null,"*","PORT_16_COUNT",port_count[16]);
	     uvm_config_db #(int)::set(null,"*","PORT_17_COUNT",port_count[17]);
	     uvm_config_db #(int)::set(null,"*","PORT_18_COUNT",port_count[18]);
	     uvm_config_db #(int)::set(null,"*","PORT_19_COUNT",port_count[19]);
	     uvm_config_db #(int)::set(null,"*","PORT_20_COUNT",port_count[20]);
	     uvm_config_db #(int)::set(null,"*","PORT_21_COUNT",port_count[21]);
	     uvm_config_db #(int)::set(null,"*","PORT_22_COUNT",port_count[22]);
	     uvm_config_db #(int)::set(null,"*","PORT_23_COUNT",port_count[23]);
       `endif
       `ifdef TB_CONFIG_3
       uvm_config_db #(int)::set(null,"*","PORT_24_COUNT",port_count[24]);
	     uvm_config_db #(int)::set(null,"*","PORT_25_COUNT",port_count[25]);
	     uvm_config_db #(int)::set(null,"*","PORT_26_COUNT",port_count[26]);
	     uvm_config_db #(int)::set(null,"*","PORT_27_COUNT",port_count[27]);
	     uvm_config_db #(int)::set(null,"*","PORT_28_COUNT",port_count[28]);
	     uvm_config_db #(int)::set(null,"*","PORT_29_COUNT",port_count[29]);
	     uvm_config_db #(int)::set(null,"*","PORT_30_COUNT",port_count[30]);
	     uvm_config_db #(int)::set(null,"*","PORT_31_COUNT",port_count[31]);
       `endif
       `ifdef TB_CONFIG_4
       uvm_config_db #(int)::set(null,"*","PORT_24_COUNT",port_count[24]);
       uvm_config_db #(int)::set(null,"*","PORT_25_COUNT",port_count[25]);
       uvm_config_db #(int)::set(null,"*","PORT_26_COUNT",port_count[26]);
       uvm_config_db #(int)::set(null,"*","PORT_27_COUNT",port_count[27]);
       uvm_config_db #(int)::set(null,"*","PORT_28_COUNT",port_count[28]);
       uvm_config_db #(int)::set(null,"*","PORT_29_COUNT",port_count[29]);
       uvm_config_db #(int)::set(null,"*","PORT_30_COUNT",port_count[30]);
       uvm_config_db #(int)::set(null,"*","PORT_31_COUNT",port_count[31]);
       uvm_config_db #(int)::set(null,"*","PORT_32_COUNT",port_count[32]);
       uvm_config_db #(int)::set(null,"*","PORT_33_COUNT",port_count[33]);
       uvm_config_db #(int)::set(null,"*","PORT_34_COUNT",port_count[34]);
       uvm_config_db #(int)::set(null,"*","PORT_35_COUNT",port_count[35]);
       uvm_config_db #(int)::set(null,"*","PORT_36_COUNT",port_count[36]);
       uvm_config_db #(int)::set(null,"*","PORT_37_COUNT",port_count[37]);
       uvm_config_db #(int)::set(null,"*","PORT_38_COUNT",port_count[38]);
       uvm_config_db #(int)::set(null,"*","PORT_39_COUNT",port_count[39]);
       uvm_config_db #(int)::set(null,"*","PORT_40_COUNT",port_count[40]);
       uvm_config_db #(int)::set(null,"*","PORT_41_COUNT",port_count[41]);
       uvm_config_db #(int)::set(null,"*","PORT_42_COUNT",port_count[42]);
       uvm_config_db #(int)::set(null,"*","PORT_43_COUNT",port_count[43]);
       uvm_config_db #(int)::set(null,"*","PORT_44_COUNT",port_count[44]);
       uvm_config_db #(int)::set(null,"*","PORT_45_COUNT",port_count[45]);
       uvm_config_db #(int)::set(null,"*","PORT_46_COUNT",port_count[46]);
       uvm_config_db #(int)::set(null,"*","PORT_47_COUNT",port_count[47]);
       uvm_config_db #(int)::set(null,"*","PORT_48_COUNT",port_count[48]);
       uvm_config_db #(int)::set(null,"*","PORT_49_COUNT",port_count[49]);
       uvm_config_db #(int)::set(null,"*","PORT_50_COUNT",port_count[50]);
       uvm_config_db #(int)::set(null,"*","PORT_51_COUNT",port_count[51]);
       uvm_config_db #(int)::set(null,"*","PORT_52_COUNT",port_count[52]);
       uvm_config_db #(int)::set(null,"*","PORT_53_COUNT",port_count[53]);
       uvm_config_db #(int)::set(null,"*","PORT_54_COUNT",port_count[54]);
       uvm_config_db #(int)::set(null,"*","PORT_55_COUNT",port_count[55]);
       uvm_config_db #(int)::set(null,"*","PORT_56_COUNT",port_count[56]);
       uvm_config_db #(int)::set(null,"*","PORT_57_COUNT",port_count[57]);
       uvm_config_db #(int)::set(null,"*","PORT_58_COUNT",port_count[58]);
       uvm_config_db #(int)::set(null,"*","PORT_59_COUNT",port_count[59]);
       uvm_config_db #(int)::set(null,"*","PORT_60_COUNT",port_count[60]);
       uvm_config_db #(int)::set(null,"*","PORT_61_COUNT",port_count[61]);
       uvm_config_db #(int)::set(null,"*","PORT_62_COUNT",port_count[62]);
       uvm_config_db #(int)::set(null,"*","PORT_63_COUNT",port_count[63]);
       uvm_config_db #(int)::set(null,"*","PORT_64_COUNT",port_count[64]);
       uvm_config_db #(int)::set(null,"*","PORT_65_COUNT",port_count[65]);
       uvm_config_db #(int)::set(null,"*","PORT_66_COUNT",port_count[66]);
       uvm_config_db #(int)::set(null,"*","PORT_67_COUNT",port_count[67]);
       uvm_config_db #(int)::set(null,"*","PORT_68_COUNT",port_count[68]);
       uvm_config_db #(int)::set(null,"*","PORT_69_COUNT",port_count[69]);
       uvm_config_db #(int)::set(null,"*","PORT_70_COUNT",port_count[70]);
       uvm_config_db #(int)::set(null,"*","PORT_71_COUNT",port_count[71]);
       uvm_config_db #(int)::set(null,"*","PORT_72_COUNT",port_count[72]);
       uvm_config_db #(int)::set(null,"*","PORT_73_COUNT",port_count[73]);
       uvm_config_db #(int)::set(null,"*","PORT_74_COUNT",port_count[74]);
       uvm_config_db #(int)::set(null,"*","PORT_75_COUNT",port_count[75]);
       uvm_config_db #(int)::set(null,"*","PORT_76_COUNT",port_count[76]);
       uvm_config_db #(int)::set(null,"*","PORT_77_COUNT",port_count[77]);
       uvm_config_db #(int)::set(null,"*","PORT_78_COUNT",port_count[78]);
       uvm_config_db #(int)::set(null,"*","PORT_79_COUNT",port_count[79]);
       uvm_config_db #(int)::set(null,"*","PORT_80_COUNT",port_count[80]);
       uvm_config_db #(int)::set(null,"*","PORT_81_COUNT",port_count[81]);
       uvm_config_db #(int)::set(null,"*","PORT_82_COUNT",port_count[82]);
       uvm_config_db #(int)::set(null,"*","PORT_83_COUNT",port_count[83]);
       uvm_config_db #(int)::set(null,"*","PORT_84_COUNT",port_count[84]);
       uvm_config_db #(int)::set(null,"*","PORT_85_COUNT",port_count[85]);
       uvm_config_db #(int)::set(null,"*","PORT_86_COUNT",port_count[86]);
       uvm_config_db #(int)::set(null,"*","PORT_87_COUNT",port_count[87]);
       uvm_config_db #(int)::set(null,"*","PORT_88_COUNT",port_count[88]);
       uvm_config_db #(int)::set(null,"*","PORT_89_COUNT",port_count[89]);
       uvm_config_db #(int)::set(null,"*","PORT_90_COUNT",port_count[90]);
       uvm_config_db #(int)::set(null,"*","PORT_91_COUNT",port_count[91]);
       uvm_config_db #(int)::set(null,"*","PORT_92_COUNT",port_count[92]);
       uvm_config_db #(int)::set(null,"*","PORT_93_COUNT",port_count[93]);
       uvm_config_db #(int)::set(null,"*","PORT_94_COUNT",port_count[94]);
       uvm_config_db #(int)::set(null,"*","PORT_95_COUNT",port_count[95]);
       uvm_config_db #(int)::set(null,"*","PORT_96_COUNT",port_count[96]);
       uvm_config_db #(int)::set(null,"*","PORT_97_COUNT",port_count[97]);
       uvm_config_db #(int)::set(null,"*","PORT_98_COUNT",port_count[98]);
       uvm_config_db #(int)::set(null,"*","PORT_99_COUNT",port_count[99]);
       uvm_config_db #(int)::set(null,"*","PORT_100_COUNT",port_count[100]);
       uvm_config_db #(int)::set(null,"*","PORT_101_COUNT",port_count[101]);
       uvm_config_db #(int)::set(null,"*","PORT_102_COUNT",port_count[102]);
       uvm_config_db #(int)::set(null,"*","PORT_103_COUNT",port_count[103]);
       uvm_config_db #(int)::set(null,"*","PORT_104_COUNT",port_count[104]);
       uvm_config_db #(int)::set(null,"*","PORT_105_COUNT",port_count[105]);
       uvm_config_db #(int)::set(null,"*","PORT_106_COUNT",port_count[106]);
       uvm_config_db #(int)::set(null,"*","PORT_107_COUNT",port_count[107]);
       uvm_config_db #(int)::set(null,"*","PORT_108_COUNT",port_count[108]);
       uvm_config_db #(int)::set(null,"*","PORT_109_COUNT",port_count[109]);
       uvm_config_db #(int)::set(null,"*","PORT_110_COUNT",port_count[110]);
       uvm_config_db #(int)::set(null,"*","PORT_111_COUNT",port_count[111]);
       uvm_config_db #(int)::set(null,"*","PORT_112_COUNT",port_count[112]);
       uvm_config_db #(int)::set(null,"*","PORT_113_COUNT",port_count[113]);
       uvm_config_db #(int)::set(null,"*","PORT_114_COUNT",port_count[114]);
       uvm_config_db #(int)::set(null,"*","PORT_115_COUNT",port_count[115]);
       uvm_config_db #(int)::set(null,"*","PORT_116_COUNT",port_count[116]);
       uvm_config_db #(int)::set(null,"*","PORT_117_COUNT",port_count[117]);
       uvm_config_db #(int)::set(null,"*","PORT_118_COUNT",port_count[118]);
       uvm_config_db #(int)::set(null,"*","PORT_119_COUNT",port_count[119]);
       uvm_config_db #(int)::set(null,"*","PORT_120_COUNT",port_count[120]);
       uvm_config_db #(int)::set(null,"*","PORT_121_COUNT",port_count[121]);
       uvm_config_db #(int)::set(null,"*","PORT_122_COUNT",port_count[122]);
       uvm_config_db #(int)::set(null,"*","PORT_123_COUNT",port_count[123]);
       uvm_config_db #(int)::set(null,"*","PORT_124_COUNT",port_count[124]);
       uvm_config_db #(int)::set(null,"*","PORT_125_COUNT",port_count[125]);
       uvm_config_db #(int)::set(null,"*","PORT_126_COUNT",port_count[126]);
       uvm_config_db #(int)::set(null,"*","PORT_127_COUNT",port_count[127]);
       uvm_config_db #(int)::set(null,"*","PORT_128_COUNT",port_count[128]);
       uvm_config_db #(int)::set(null,"*","PORT_129_COUNT",port_count[129]);
       uvm_config_db #(int)::set(null,"*","PORT_130_COUNT",port_count[130]);
       uvm_config_db #(int)::set(null,"*","PORT_131_COUNT",port_count[131]);
       uvm_config_db #(int)::set(null,"*","PORT_132_COUNT",port_count[132]);
       uvm_config_db #(int)::set(null,"*","PORT_133_COUNT",port_count[133]);
       uvm_config_db #(int)::set(null,"*","PORT_134_COUNT",port_count[134]);
       uvm_config_db #(int)::set(null,"*","PORT_135_COUNT",port_count[135]);
       uvm_config_db #(int)::set(null,"*","PORT_136_COUNT",port_count[136]);
       uvm_config_db #(int)::set(null,"*","PORT_137_COUNT",port_count[137]);
       uvm_config_db #(int)::set(null,"*","PORT_138_COUNT",port_count[138]);
       uvm_config_db #(int)::set(null,"*","PORT_139_COUNT",port_count[139]);
       uvm_config_db #(int)::set(null,"*","PORT_140_COUNT",port_count[140]);
       uvm_config_db #(int)::set(null,"*","PORT_141_COUNT",port_count[141]);
       uvm_config_db #(int)::set(null,"*","PORT_142_COUNT",port_count[142]);
       uvm_config_db #(int)::set(null,"*","PORT_143_COUNT",port_count[143]);
       uvm_config_db #(int)::set(null,"*","PORT_144_COUNT",port_count[144]);
       uvm_config_db #(int)::set(null,"*","PORT_145_COUNT",port_count[145]);
       uvm_config_db #(int)::set(null,"*","PORT_146_COUNT",port_count[146]);
       uvm_config_db #(int)::set(null,"*","PORT_147_COUNT",port_count[147]);
       uvm_config_db #(int)::set(null,"*","PORT_148_COUNT",port_count[148]);
       uvm_config_db #(int)::set(null,"*","PORT_149_COUNT",port_count[149]);
       uvm_config_db #(int)::set(null,"*","PORT_150_COUNT",port_count[150]);
       uvm_config_db #(int)::set(null,"*","PORT_151_COUNT",port_count[151]);
       uvm_config_db #(int)::set(null,"*","PORT_152_COUNT",port_count[152]);
       uvm_config_db #(int)::set(null,"*","PORT_153_COUNT",port_count[153]);
       uvm_config_db #(int)::set(null,"*","PORT_154_COUNT",port_count[154]);
       uvm_config_db #(int)::set(null,"*","PORT_155_COUNT",port_count[155]);
       uvm_config_db #(int)::set(null,"*","PORT_156_COUNT",port_count[156]);
       uvm_config_db #(int)::set(null,"*","PORT_157_COUNT",port_count[157]);
       uvm_config_db #(int)::set(null,"*","PORT_158_COUNT",port_count[158]);
       uvm_config_db #(int)::set(null,"*","PORT_159_COUNT",port_count[159]);
       uvm_config_db #(int)::set(null,"*","PORT_160_COUNT",port_count[160]);
       uvm_config_db #(int)::set(null,"*","PORT_161_COUNT",port_count[161]);
       uvm_config_db #(int)::set(null,"*","PORT_162_COUNT",port_count[162]);
       uvm_config_db #(int)::set(null,"*","PORT_163_COUNT",port_count[163]);
       uvm_config_db #(int)::set(null,"*","PORT_164_COUNT",port_count[164]);
       uvm_config_db #(int)::set(null,"*","PORT_165_COUNT",port_count[165]);
       uvm_config_db #(int)::set(null,"*","PORT_166_COUNT",port_count[166]);
       uvm_config_db #(int)::set(null,"*","PORT_167_COUNT",port_count[167]);
       uvm_config_db #(int)::set(null,"*","PORT_168_COUNT",port_count[168]);
       uvm_config_db #(int)::set(null,"*","PORT_169_COUNT",port_count[169]);
       uvm_config_db #(int)::set(null,"*","PORT_170_COUNT",port_count[170]);
       uvm_config_db #(int)::set(null,"*","PORT_171_COUNT",port_count[171]);
       uvm_config_db #(int)::set(null,"*","PORT_172_COUNT",port_count[172]);
       uvm_config_db #(int)::set(null,"*","PORT_173_COUNT",port_count[173]);
       uvm_config_db #(int)::set(null,"*","PORT_174_COUNT",port_count[174]);
       uvm_config_db #(int)::set(null,"*","PORT_175_COUNT",port_count[175]);
       uvm_config_db #(int)::set(null,"*","PORT_176_COUNT",port_count[176]);
       uvm_config_db #(int)::set(null,"*","PORT_177_COUNT",port_count[177]);
       uvm_config_db #(int)::set(null,"*","PORT_178_COUNT",port_count[178]);
       uvm_config_db #(int)::set(null,"*","PORT_179_COUNT",port_count[179]);
       uvm_config_db #(int)::set(null,"*","PORT_180_COUNT",port_count[180]);
       uvm_config_db #(int)::set(null,"*","PORT_181_COUNT",port_count[181]);
       uvm_config_db #(int)::set(null,"*","PORT_182_COUNT",port_count[182]);
       uvm_config_db #(int)::set(null,"*","PORT_183_COUNT",port_count[183]);
       uvm_config_db #(int)::set(null,"*","PORT_184_COUNT",port_count[184]);
       uvm_config_db #(int)::set(null,"*","PORT_185_COUNT",port_count[185]);
       uvm_config_db #(int)::set(null,"*","PORT_186_COUNT",port_count[186]);
       uvm_config_db #(int)::set(null,"*","PORT_187_COUNT",port_count[187]);
       uvm_config_db #(int)::set(null,"*","PORT_188_COUNT",port_count[188]);
       uvm_config_db #(int)::set(null,"*","PORT_189_COUNT",port_count[189]);
       uvm_config_db #(int)::set(null,"*","PORT_190_COUNT",port_count[190]);
       uvm_config_db #(int)::set(null,"*","PORT_191_COUNT",port_count[191]);
       uvm_config_db #(int)::set(null,"*","PORT_192_COUNT",port_count[192]);
       uvm_config_db #(int)::set(null,"*","PORT_193_COUNT",port_count[193]);
       uvm_config_db #(int)::set(null,"*","PORT_194_COUNT",port_count[194]);
       uvm_config_db #(int)::set(null,"*","PORT_195_COUNT",port_count[195]);
       uvm_config_db #(int)::set(null,"*","PORT_196_COUNT",port_count[196]);
       uvm_config_db #(int)::set(null,"*","PORT_197_COUNT",port_count[197]);
       uvm_config_db #(int)::set(null,"*","PORT_198_COUNT",port_count[198]);
       uvm_config_db #(int)::set(null,"*","PORT_199_COUNT",port_count[199]);
       uvm_config_db #(int)::set(null,"*","PORT_200_COUNT",port_count[200]);
       uvm_config_db #(int)::set(null,"*","PORT_201_COUNT",port_count[201]);
       uvm_config_db #(int)::set(null,"*","PORT_202_COUNT",port_count[202]);
       uvm_config_db #(int)::set(null,"*","PORT_203_COUNT",port_count[203]);
       uvm_config_db #(int)::set(null,"*","PORT_204_COUNT",port_count[204]);
       uvm_config_db #(int)::set(null,"*","PORT_205_COUNT",port_count[205]);
       uvm_config_db #(int)::set(null,"*","PORT_206_COUNT",port_count[206]);
       uvm_config_db #(int)::set(null,"*","PORT_207_COUNT",port_count[207]);
       uvm_config_db #(int)::set(null,"*","PORT_208_COUNT",port_count[208]);
       uvm_config_db #(int)::set(null,"*","PORT_209_COUNT",port_count[209]);
       uvm_config_db #(int)::set(null,"*","PORT_210_COUNT",port_count[210]);
       uvm_config_db #(int)::set(null,"*","PORT_211_COUNT",port_count[211]);
       uvm_config_db #(int)::set(null,"*","PORT_212_COUNT",port_count[212]);
       uvm_config_db #(int)::set(null,"*","PORT_213_COUNT",port_count[213]);
       uvm_config_db #(int)::set(null,"*","PORT_214_COUNT",port_count[214]);
       uvm_config_db #(int)::set(null,"*","PORT_215_COUNT",port_count[215]);
       uvm_config_db #(int)::set(null,"*","PORT_216_COUNT",port_count[216]);
       uvm_config_db #(int)::set(null,"*","PORT_217_COUNT",port_count[217]);
       uvm_config_db #(int)::set(null,"*","PORT_218_COUNT",port_count[218]);
       uvm_config_db #(int)::set(null,"*","PORT_219_COUNT",port_count[219]);
       uvm_config_db #(int)::set(null,"*","PORT_220_COUNT",port_count[220]);
       uvm_config_db #(int)::set(null,"*","PORT_221_COUNT",port_count[221]);
       uvm_config_db #(int)::set(null,"*","PORT_222_COUNT",port_count[222]);
       uvm_config_db #(int)::set(null,"*","PORT_223_COUNT",port_count[223]);
       uvm_config_db #(int)::set(null,"*","PORT_224_COUNT",port_count[224]);
       uvm_config_db #(int)::set(null,"*","PORT_225_COUNT",port_count[225]);
       uvm_config_db #(int)::set(null,"*","PORT_226_COUNT",port_count[226]);
       uvm_config_db #(int)::set(null,"*","PORT_227_COUNT",port_count[227]);
       uvm_config_db #(int)::set(null,"*","PORT_228_COUNT",port_count[228]);
       uvm_config_db #(int)::set(null,"*","PORT_229_COUNT",port_count[229]);
       uvm_config_db #(int)::set(null,"*","PORT_230_COUNT",port_count[230]);
       uvm_config_db #(int)::set(null,"*","PORT_231_COUNT",port_count[231]);
       uvm_config_db #(int)::set(null,"*","PORT_232_COUNT",port_count[232]);
       uvm_config_db #(int)::set(null,"*","PORT_233_COUNT",port_count[233]);
       uvm_config_db #(int)::set(null,"*","PORT_234_COUNT",port_count[234]);
       uvm_config_db #(int)::set(null,"*","PORT_235_COUNT",port_count[235]);
       uvm_config_db #(int)::set(null,"*","PORT_236_COUNT",port_count[236]);
       uvm_config_db #(int)::set(null,"*","PORT_237_COUNT",port_count[237]);
       uvm_config_db #(int)::set(null,"*","PORT_238_COUNT",port_count[238]);
       uvm_config_db #(int)::set(null,"*","PORT_239_COUNT",port_count[239]);
       uvm_config_db #(int)::set(null,"*","PORT_240_COUNT",port_count[240]);
       uvm_config_db #(int)::set(null,"*","PORT_241_COUNT",port_count[241]);
       uvm_config_db #(int)::set(null,"*","PORT_242_COUNT",port_count[242]);
       uvm_config_db #(int)::set(null,"*","PORT_243_COUNT",port_count[243]);
       uvm_config_db #(int)::set(null,"*","PORT_244_COUNT",port_count[244]);
       uvm_config_db #(int)::set(null,"*","PORT_245_COUNT",port_count[245]);
       uvm_config_db #(int)::set(null,"*","PORT_246_COUNT",port_count[246]);
       uvm_config_db #(int)::set(null,"*","PORT_247_COUNT",port_count[247]);
       uvm_config_db #(int)::set(null,"*","PORT_248_COUNT",port_count[248]);
       uvm_config_db #(int)::set(null,"*","PORT_249_COUNT",port_count[249]);
       uvm_config_db #(int)::set(null,"*","PORT_250_COUNT",port_count[250]);
       uvm_config_db #(int)::set(null,"*","PORT_251_COUNT",port_count[251]);
       uvm_config_db #(int)::set(null,"*","PORT_252_COUNT",port_count[252]);
       uvm_config_db #(int)::set(null,"*","PORT_253_COUNT",port_count[253]);
       uvm_config_db #(int)::set(null,"*","PORT_254_COUNT",port_count[254]);
       uvm_config_db #(int)::set(null,"*","PORT_255_COUNT",port_count[255]);
       uvm_config_db #(int)::set(null,"*","PORT_256_COUNT",port_count[256]);
       uvm_config_db #(int)::set(null,"*","PORT_257_COUNT",port_count[257]);
       uvm_config_db #(int)::set(null,"*","PORT_258_COUNT",port_count[258]);
       uvm_config_db #(int)::set(null,"*","PORT_259_COUNT",port_count[259]);
       uvm_config_db #(int)::set(null,"*","PORT_260_COUNT",port_count[260]);
       uvm_config_db #(int)::set(null,"*","PORT_261_COUNT",port_count[261]);
       uvm_config_db #(int)::set(null,"*","PORT_262_COUNT",port_count[262]);
       uvm_config_db #(int)::set(null,"*","PORT_263_COUNT",port_count[263]);
       uvm_config_db #(int)::set(null,"*","PORT_264_COUNT",port_count[264]);
       uvm_config_db #(int)::set(null,"*","PORT_265_COUNT",port_count[265]);
       uvm_config_db #(int)::set(null,"*","PORT_266_COUNT",port_count[266]);
       uvm_config_db #(int)::set(null,"*","PORT_267_COUNT",port_count[267]);
       uvm_config_db #(int)::set(null,"*","PORT_268_COUNT",port_count[268]);
       uvm_config_db #(int)::set(null,"*","PORT_269_COUNT",port_count[269]);
       uvm_config_db #(int)::set(null,"*","PORT_270_COUNT",port_count[270]);
       uvm_config_db #(int)::set(null,"*","PORT_271_COUNT",port_count[271]);
       uvm_config_db #(int)::set(null,"*","PORT_272_COUNT",port_count[272]);
       uvm_config_db #(int)::set(null,"*","PORT_273_COUNT",port_count[273]);
       uvm_config_db #(int)::set(null,"*","PORT_274_COUNT",port_count[274]);
       uvm_config_db #(int)::set(null,"*","PORT_275_COUNT",port_count[275]);
       uvm_config_db #(int)::set(null,"*","PORT_276_COUNT",port_count[276]);
       uvm_config_db #(int)::set(null,"*","PORT_277_COUNT",port_count[277]);
       uvm_config_db #(int)::set(null,"*","PORT_278_COUNT",port_count[278]);
       uvm_config_db #(int)::set(null,"*","PORT_279_COUNT",port_count[279]);
       uvm_config_db #(int)::set(null,"*","PORT_280_COUNT",port_count[280]);
       uvm_config_db #(int)::set(null,"*","PORT_281_COUNT",port_count[281]);
       uvm_config_db #(int)::set(null,"*","PORT_282_COUNT",port_count[282]);
       uvm_config_db #(int)::set(null,"*","PORT_283_COUNT",port_count[283]);
       uvm_config_db #(int)::set(null,"*","PORT_284_COUNT",port_count[284]);
       uvm_config_db #(int)::set(null,"*","PORT_285_COUNT",port_count[285]);
       uvm_config_db #(int)::set(null,"*","PORT_286_COUNT",port_count[286]);
       uvm_config_db #(int)::set(null,"*","PORT_287_COUNT",port_count[287]);
       uvm_config_db #(int)::set(null,"*","PORT_288_COUNT",port_count[288]);
       uvm_config_db #(int)::set(null,"*","PORT_289_COUNT",port_count[289]);
       uvm_config_db #(int)::set(null,"*","PORT_290_COUNT",port_count[290]);
       uvm_config_db #(int)::set(null,"*","PORT_291_COUNT",port_count[291]);
       uvm_config_db #(int)::set(null,"*","PORT_292_COUNT",port_count[292]);
       uvm_config_db #(int)::set(null,"*","PORT_293_COUNT",port_count[293]);
       uvm_config_db #(int)::set(null,"*","PORT_294_COUNT",port_count[294]);
       uvm_config_db #(int)::set(null,"*","PORT_295_COUNT",port_count[295]);
       uvm_config_db #(int)::set(null,"*","PORT_296_COUNT",port_count[296]);
       uvm_config_db #(int)::set(null,"*","PORT_297_COUNT",port_count[297]);
       uvm_config_db #(int)::set(null,"*","PORT_298_COUNT",port_count[298]);
       uvm_config_db #(int)::set(null,"*","PORT_299_COUNT",port_count[299]);
       uvm_config_db #(int)::set(null,"*","PORT_300_COUNT",port_count[300]);
       uvm_config_db #(int)::set(null,"*","PORT_301_COUNT",port_count[301]);
       uvm_config_db #(int)::set(null,"*","PORT_302_COUNT",port_count[302]);
       uvm_config_db #(int)::set(null,"*","PORT_303_COUNT",port_count[303]);
       uvm_config_db #(int)::set(null,"*","PORT_304_COUNT",port_count[304]);
       uvm_config_db #(int)::set(null,"*","PORT_305_COUNT",port_count[305]);
       uvm_config_db #(int)::set(null,"*","PORT_306_COUNT",port_count[306]);
       uvm_config_db #(int)::set(null,"*","PORT_307_COUNT",port_count[307]);
       uvm_config_db #(int)::set(null,"*","PORT_308_COUNT",port_count[308]);
       uvm_config_db #(int)::set(null,"*","PORT_309_COUNT",port_count[309]);
       uvm_config_db #(int)::set(null,"*","PORT_310_COUNT",port_count[310]);
       uvm_config_db #(int)::set(null,"*","PORT_311_COUNT",port_count[311]);
       uvm_config_db #(int)::set(null,"*","PORT_312_COUNT",port_count[312]);
       uvm_config_db #(int)::set(null,"*","PORT_313_COUNT",port_count[313]);
       uvm_config_db #(int)::set(null,"*","PORT_314_COUNT",port_count[314]);
       uvm_config_db #(int)::set(null,"*","PORT_315_COUNT",port_count[315]);
       uvm_config_db #(int)::set(null,"*","PORT_316_COUNT",port_count[316]);
       uvm_config_db #(int)::set(null,"*","PORT_317_COUNT",port_count[317]);
       uvm_config_db #(int)::set(null,"*","PORT_318_COUNT",port_count[318]);
       uvm_config_db #(int)::set(null,"*","PORT_319_COUNT",port_count[319]);
       uvm_config_db #(int)::set(null,"*","PORT_320_COUNT",port_count[320]);
       uvm_config_db #(int)::set(null,"*","PORT_321_COUNT",port_count[321]);
       uvm_config_db #(int)::set(null,"*","PORT_322_COUNT",port_count[322]);
       uvm_config_db #(int)::set(null,"*","PORT_323_COUNT",port_count[323]);
       uvm_config_db #(int)::set(null,"*","PORT_324_COUNT",port_count[324]);
       uvm_config_db #(int)::set(null,"*","PORT_325_COUNT",port_count[325]);
       uvm_config_db #(int)::set(null,"*","PORT_326_COUNT",port_count[326]);
       uvm_config_db #(int)::set(null,"*","PORT_327_COUNT",port_count[327]);
       uvm_config_db #(int)::set(null,"*","PORT_328_COUNT",port_count[328]);
       uvm_config_db #(int)::set(null,"*","PORT_329_COUNT",port_count[329]);
       uvm_config_db #(int)::set(null,"*","PORT_330_COUNT",port_count[330]);
       uvm_config_db #(int)::set(null,"*","PORT_331_COUNT",port_count[331]);
       uvm_config_db #(int)::set(null,"*","PORT_332_COUNT",port_count[332]);
       uvm_config_db #(int)::set(null,"*","PORT_333_COUNT",port_count[333]);
       uvm_config_db #(int)::set(null,"*","PORT_334_COUNT",port_count[334]);
       uvm_config_db #(int)::set(null,"*","PORT_335_COUNT",port_count[335]);
       uvm_config_db #(int)::set(null,"*","PORT_336_COUNT",port_count[336]);
       uvm_config_db #(int)::set(null,"*","PORT_337_COUNT",port_count[337]);
       uvm_config_db #(int)::set(null,"*","PORT_338_COUNT",port_count[338]);
       uvm_config_db #(int)::set(null,"*","PORT_339_COUNT",port_count[339]);
       uvm_config_db #(int)::set(null,"*","PORT_340_COUNT",port_count[340]);
       uvm_config_db #(int)::set(null,"*","PORT_341_COUNT",port_count[341]);
       uvm_config_db #(int)::set(null,"*","PORT_342_COUNT",port_count[342]);
       uvm_config_db #(int)::set(null,"*","PORT_343_COUNT",port_count[343]);
       uvm_config_db #(int)::set(null,"*","PORT_344_COUNT",port_count[344]);
       uvm_config_db #(int)::set(null,"*","PORT_345_COUNT",port_count[345]);
       uvm_config_db #(int)::set(null,"*","PORT_346_COUNT",port_count[346]);
       uvm_config_db #(int)::set(null,"*","PORT_347_COUNT",port_count[347]);
       uvm_config_db #(int)::set(null,"*","PORT_348_COUNT",port_count[348]);
       uvm_config_db #(int)::set(null,"*","PORT_349_COUNT",port_count[349]);
       uvm_config_db #(int)::set(null,"*","PORT_350_COUNT",port_count[350]);
       uvm_config_db #(int)::set(null,"*","PORT_351_COUNT",port_count[351]);
       uvm_config_db #(int)::set(null,"*","PORT_352_COUNT",port_count[352]);
       uvm_config_db #(int)::set(null,"*","PORT_353_COUNT",port_count[353]);
       uvm_config_db #(int)::set(null,"*","PORT_354_COUNT",port_count[354]);
       uvm_config_db #(int)::set(null,"*","PORT_355_COUNT",port_count[355]);
       uvm_config_db #(int)::set(null,"*","PORT_356_COUNT",port_count[356]);
       uvm_config_db #(int)::set(null,"*","PORT_357_COUNT",port_count[357]);
       uvm_config_db #(int)::set(null,"*","PORT_358_COUNT",port_count[358]);
       uvm_config_db #(int)::set(null,"*","PORT_359_COUNT",port_count[359]);
       uvm_config_db #(int)::set(null,"*","PORT_360_COUNT",port_count[360]);
       uvm_config_db #(int)::set(null,"*","PORT_361_COUNT",port_count[361]);
       uvm_config_db #(int)::set(null,"*","PORT_362_COUNT",port_count[362]);
       uvm_config_db #(int)::set(null,"*","PORT_363_COUNT",port_count[363]);
       uvm_config_db #(int)::set(null,"*","PORT_364_COUNT",port_count[364]);
       uvm_config_db #(int)::set(null,"*","PORT_365_COUNT",port_count[365]);
       uvm_config_db #(int)::set(null,"*","PORT_366_COUNT",port_count[366]);
       uvm_config_db #(int)::set(null,"*","PORT_367_COUNT",port_count[367]);
       uvm_config_db #(int)::set(null,"*","PORT_368_COUNT",port_count[368]);
       uvm_config_db #(int)::set(null,"*","PORT_369_COUNT",port_count[369]);
       uvm_config_db #(int)::set(null,"*","PORT_370_COUNT",port_count[370]);
       uvm_config_db #(int)::set(null,"*","PORT_371_COUNT",port_count[371]);
       uvm_config_db #(int)::set(null,"*","PORT_372_COUNT",port_count[372]);
       uvm_config_db #(int)::set(null,"*","PORT_373_COUNT",port_count[373]);
       uvm_config_db #(int)::set(null,"*","PORT_374_COUNT",port_count[374]);
       uvm_config_db #(int)::set(null,"*","PORT_375_COUNT",port_count[375]);
       uvm_config_db #(int)::set(null,"*","PORT_376_COUNT",port_count[376]);
       uvm_config_db #(int)::set(null,"*","PORT_377_COUNT",port_count[377]);
       uvm_config_db #(int)::set(null,"*","PORT_378_COUNT",port_count[378]);
       uvm_config_db #(int)::set(null,"*","PORT_379_COUNT",port_count[379]);
       uvm_config_db #(int)::set(null,"*","PORT_380_COUNT",port_count[380]);
       uvm_config_db #(int)::set(null,"*","PORT_381_COUNT",port_count[381]);
       uvm_config_db #(int)::set(null,"*","PORT_382_COUNT",port_count[382]);
       uvm_config_db #(int)::set(null,"*","PORT_383_COUNT",port_count[383]);
       uvm_config_db #(int)::set(null,"*","PORT_384_COUNT",port_count[384]);
       uvm_config_db #(int)::set(null,"*","PORT_385_COUNT",port_count[385]);
       uvm_config_db #(int)::set(null,"*","PORT_386_COUNT",port_count[386]);
       uvm_config_db #(int)::set(null,"*","PORT_387_COUNT",port_count[387]);
       uvm_config_db #(int)::set(null,"*","PORT_388_COUNT",port_count[388]);
       uvm_config_db #(int)::set(null,"*","PORT_389_COUNT",port_count[389]);
       uvm_config_db #(int)::set(null,"*","PORT_390_COUNT",port_count[390]);
       uvm_config_db #(int)::set(null,"*","PORT_391_COUNT",port_count[391]);
       uvm_config_db #(int)::set(null,"*","PORT_392_COUNT",port_count[392]);
       uvm_config_db #(int)::set(null,"*","PORT_393_COUNT",port_count[393]);
       uvm_config_db #(int)::set(null,"*","PORT_394_COUNT",port_count[394]);
       uvm_config_db #(int)::set(null,"*","PORT_395_COUNT",port_count[395]);
       uvm_config_db #(int)::set(null,"*","PORT_396_COUNT",port_count[396]);
       uvm_config_db #(int)::set(null,"*","PORT_397_COUNT",port_count[397]);
       uvm_config_db #(int)::set(null,"*","PORT_398_COUNT",port_count[398]);
       uvm_config_db #(int)::set(null,"*","PORT_399_COUNT",port_count[399]);
       uvm_config_db #(int)::set(null,"*","PORT_400_COUNT",port_count[400]);
       uvm_config_db #(int)::set(null,"*","PORT_401_COUNT",port_count[401]);
       uvm_config_db #(int)::set(null,"*","PORT_402_COUNT",port_count[402]);
       uvm_config_db #(int)::set(null,"*","PORT_403_COUNT",port_count[403]);
       uvm_config_db #(int)::set(null,"*","PORT_404_COUNT",port_count[404]);
       uvm_config_db #(int)::set(null,"*","PORT_405_COUNT",port_count[405]);
       uvm_config_db #(int)::set(null,"*","PORT_406_COUNT",port_count[406]);
       uvm_config_db #(int)::set(null,"*","PORT_407_COUNT",port_count[407]);
       uvm_config_db #(int)::set(null,"*","PORT_408_COUNT",port_count[408]);
       uvm_config_db #(int)::set(null,"*","PORT_409_COUNT",port_count[409]);
       uvm_config_db #(int)::set(null,"*","PORT_410_COUNT",port_count[410]);
       uvm_config_db #(int)::set(null,"*","PORT_411_COUNT",port_count[411]);
       uvm_config_db #(int)::set(null,"*","PORT_412_COUNT",port_count[412]);
       uvm_config_db #(int)::set(null,"*","PORT_413_COUNT",port_count[413]);
       uvm_config_db #(int)::set(null,"*","PORT_414_COUNT",port_count[414]);
       uvm_config_db #(int)::set(null,"*","PORT_415_COUNT",port_count[415]);
       uvm_config_db #(int)::set(null,"*","PORT_416_COUNT",port_count[416]);
       uvm_config_db #(int)::set(null,"*","PORT_417_COUNT",port_count[417]);
       uvm_config_db #(int)::set(null,"*","PORT_418_COUNT",port_count[418]);
       uvm_config_db #(int)::set(null,"*","PORT_419_COUNT",port_count[419]);
       uvm_config_db #(int)::set(null,"*","PORT_420_COUNT",port_count[420]);
       uvm_config_db #(int)::set(null,"*","PORT_421_COUNT",port_count[421]);
       uvm_config_db #(int)::set(null,"*","PORT_422_COUNT",port_count[422]);
       uvm_config_db #(int)::set(null,"*","PORT_423_COUNT",port_count[423]);
       uvm_config_db #(int)::set(null,"*","PORT_424_COUNT",port_count[424]);
       uvm_config_db #(int)::set(null,"*","PORT_425_COUNT",port_count[425]);
       uvm_config_db #(int)::set(null,"*","PORT_426_COUNT",port_count[426]);
       uvm_config_db #(int)::set(null,"*","PORT_427_COUNT",port_count[427]);
       uvm_config_db #(int)::set(null,"*","PORT_428_COUNT",port_count[428]);
       uvm_config_db #(int)::set(null,"*","PORT_429_COUNT",port_count[429]);
       uvm_config_db #(int)::set(null,"*","PORT_430_COUNT",port_count[430]);
       uvm_config_db #(int)::set(null,"*","PORT_431_COUNT",port_count[431]);
       uvm_config_db #(int)::set(null,"*","PORT_432_COUNT",port_count[432]);
       uvm_config_db #(int)::set(null,"*","PORT_433_COUNT",port_count[433]);
       uvm_config_db #(int)::set(null,"*","PORT_434_COUNT",port_count[434]);
       uvm_config_db #(int)::set(null,"*","PORT_435_COUNT",port_count[435]);
       uvm_config_db #(int)::set(null,"*","PORT_436_COUNT",port_count[436]);
       uvm_config_db #(int)::set(null,"*","PORT_437_COUNT",port_count[437]);
       uvm_config_db #(int)::set(null,"*","PORT_438_COUNT",port_count[438]);
       uvm_config_db #(int)::set(null,"*","PORT_439_COUNT",port_count[439]);
       uvm_config_db #(int)::set(null,"*","PORT_440_COUNT",port_count[440]);
       uvm_config_db #(int)::set(null,"*","PORT_441_COUNT",port_count[441]);
       uvm_config_db #(int)::set(null,"*","PORT_442_COUNT",port_count[442]);
       uvm_config_db #(int)::set(null,"*","PORT_443_COUNT",port_count[443]);
       uvm_config_db #(int)::set(null,"*","PORT_444_COUNT",port_count[444]);
       uvm_config_db #(int)::set(null,"*","PORT_445_COUNT",port_count[445]);
       uvm_config_db #(int)::set(null,"*","PORT_446_COUNT",port_count[446]);
       uvm_config_db #(int)::set(null,"*","PORT_447_COUNT",port_count[447]);
       uvm_config_db #(int)::set(null,"*","PORT_448_COUNT",port_count[448]);
       uvm_config_db #(int)::set(null,"*","PORT_449_COUNT",port_count[449]);
       uvm_config_db #(int)::set(null,"*","PORT_450_COUNT",port_count[450]);
       uvm_config_db #(int)::set(null,"*","PORT_451_COUNT",port_count[451]);
       uvm_config_db #(int)::set(null,"*","PORT_452_COUNT",port_count[452]);
       uvm_config_db #(int)::set(null,"*","PORT_453_COUNT",port_count[453]);
       uvm_config_db #(int)::set(null,"*","PORT_454_COUNT",port_count[454]);
       uvm_config_db #(int)::set(null,"*","PORT_455_COUNT",port_count[455]);
       uvm_config_db #(int)::set(null,"*","PORT_456_COUNT",port_count[456]);
       uvm_config_db #(int)::set(null,"*","PORT_457_COUNT",port_count[457]);
       uvm_config_db #(int)::set(null,"*","PORT_458_COUNT",port_count[458]);
       uvm_config_db #(int)::set(null,"*","PORT_459_COUNT",port_count[459]);
       uvm_config_db #(int)::set(null,"*","PORT_460_COUNT",port_count[460]);
       uvm_config_db #(int)::set(null,"*","PORT_461_COUNT",port_count[461]);
       uvm_config_db #(int)::set(null,"*","PORT_462_COUNT",port_count[462]);
       uvm_config_db #(int)::set(null,"*","PORT_463_COUNT",port_count[463]);
       uvm_config_db #(int)::set(null,"*","PORT_464_COUNT",port_count[464]);
       uvm_config_db #(int)::set(null,"*","PORT_465_COUNT",port_count[465]);
       uvm_config_db #(int)::set(null,"*","PORT_466_COUNT",port_count[466]);
       uvm_config_db #(int)::set(null,"*","PORT_467_COUNT",port_count[467]);
       uvm_config_db #(int)::set(null,"*","PORT_468_COUNT",port_count[468]);
       uvm_config_db #(int)::set(null,"*","PORT_469_COUNT",port_count[469]);
       uvm_config_db #(int)::set(null,"*","PORT_470_COUNT",port_count[470]);
       uvm_config_db #(int)::set(null,"*","PORT_471_COUNT",port_count[471]);
       uvm_config_db #(int)::set(null,"*","PORT_472_COUNT",port_count[472]);
       uvm_config_db #(int)::set(null,"*","PORT_473_COUNT",port_count[473]);
       uvm_config_db #(int)::set(null,"*","PORT_474_COUNT",port_count[474]);
       uvm_config_db #(int)::set(null,"*","PORT_475_COUNT",port_count[475]);
       uvm_config_db #(int)::set(null,"*","PORT_476_COUNT",port_count[476]);
       uvm_config_db #(int)::set(null,"*","PORT_477_COUNT",port_count[477]);
       uvm_config_db #(int)::set(null,"*","PORT_478_COUNT",port_count[478]);
       uvm_config_db #(int)::set(null,"*","PORT_479_COUNT",port_count[479]);
       uvm_config_db #(int)::set(null,"*","PORT_480_COUNT",port_count[480]);
       uvm_config_db #(int)::set(null,"*","PORT_481_COUNT",port_count[481]);
       uvm_config_db #(int)::set(null,"*","PORT_482_COUNT",port_count[482]);
       uvm_config_db #(int)::set(null,"*","PORT_483_COUNT",port_count[483]);
       uvm_config_db #(int)::set(null,"*","PORT_484_COUNT",port_count[484]);
       uvm_config_db #(int)::set(null,"*","PORT_485_COUNT",port_count[485]);
       uvm_config_db #(int)::set(null,"*","PORT_486_COUNT",port_count[486]);
       uvm_config_db #(int)::set(null,"*","PORT_487_COUNT",port_count[487]);
       uvm_config_db #(int)::set(null,"*","PORT_488_COUNT",port_count[488]);
       uvm_config_db #(int)::set(null,"*","PORT_489_COUNT",port_count[489]);
       uvm_config_db #(int)::set(null,"*","PORT_490_COUNT",port_count[490]);
       uvm_config_db #(int)::set(null,"*","PORT_491_COUNT",port_count[491]);
       uvm_config_db #(int)::set(null,"*","PORT_492_COUNT",port_count[492]);
       uvm_config_db #(int)::set(null,"*","PORT_493_COUNT",port_count[493]);
       uvm_config_db #(int)::set(null,"*","PORT_494_COUNT",port_count[494]);
       uvm_config_db #(int)::set(null,"*","PORT_495_COUNT",port_count[495]);
       uvm_config_db #(int)::set(null,"*","PORT_496_COUNT",port_count[496]);
       uvm_config_db #(int)::set(null,"*","PORT_497_COUNT",port_count[497]);
       uvm_config_db #(int)::set(null,"*","PORT_498_COUNT",port_count[498]);
       uvm_config_db #(int)::set(null,"*","PORT_499_COUNT",port_count[499]);
       uvm_config_db #(int)::set(null,"*","PORT_500_COUNT",port_count[500]);
       uvm_config_db #(int)::set(null,"*","PORT_501_COUNT",port_count[501]);
       uvm_config_db #(int)::set(null,"*","PORT_502_COUNT",port_count[502]);
       uvm_config_db #(int)::set(null,"*","PORT_503_COUNT",port_count[503]);
       uvm_config_db #(int)::set(null,"*","PORT_504_COUNT",port_count[504]);
       uvm_config_db #(int)::set(null,"*","PORT_505_COUNT",port_count[505]);
       uvm_config_db #(int)::set(null,"*","PORT_506_COUNT",port_count[506]);
       uvm_config_db #(int)::set(null,"*","PORT_507_COUNT",port_count[507]);
       uvm_config_db #(int)::set(null,"*","PORT_508_COUNT",port_count[508]);
       uvm_config_db #(int)::set(null,"*","PORT_509_COUNT",port_count[509]);
       uvm_config_db #(int)::set(null,"*","PORT_510_COUNT",port_count[510]);
       uvm_config_db #(int)::set(null,"*","PORT_511_COUNT",port_count[511]);
       uvm_config_db #(int)::set(null,"*","PORT_512_COUNT",port_count[512]);
       uvm_config_db #(int)::set(null,"*","PORT_513_COUNT",port_count[513]);
       uvm_config_db #(int)::set(null,"*","PORT_514_COUNT",port_count[514]);
       uvm_config_db #(int)::set(null,"*","PORT_515_COUNT",port_count[515]);
       uvm_config_db #(int)::set(null,"*","PORT_516_COUNT",port_count[516]);
       uvm_config_db #(int)::set(null,"*","PORT_517_COUNT",port_count[517]);
       uvm_config_db #(int)::set(null,"*","PORT_518_COUNT",port_count[518]);
       uvm_config_db #(int)::set(null,"*","PORT_519_COUNT",port_count[519]);
       uvm_config_db #(int)::set(null,"*","PORT_520_COUNT",port_count[520]);
       uvm_config_db #(int)::set(null,"*","PORT_521_COUNT",port_count[521]);
       uvm_config_db #(int)::set(null,"*","PORT_522_COUNT",port_count[522]);
       uvm_config_db #(int)::set(null,"*","PORT_523_COUNT",port_count[523]);
       uvm_config_db #(int)::set(null,"*","PORT_524_COUNT",port_count[524]);
       uvm_config_db #(int)::set(null,"*","PORT_525_COUNT",port_count[525]);
       uvm_config_db #(int)::set(null,"*","PORT_526_COUNT",port_count[526]);
       uvm_config_db #(int)::set(null,"*","PORT_527_COUNT",port_count[527]);
       uvm_config_db #(int)::set(null,"*","PORT_528_COUNT",port_count[528]);
       uvm_config_db #(int)::set(null,"*","PORT_529_COUNT",port_count[529]);
       uvm_config_db #(int)::set(null,"*","PORT_530_COUNT",port_count[530]);
       uvm_config_db #(int)::set(null,"*","PORT_531_COUNT",port_count[531]);
       uvm_config_db #(int)::set(null,"*","PORT_532_COUNT",port_count[532]);
       uvm_config_db #(int)::set(null,"*","PORT_533_COUNT",port_count[533]);
       uvm_config_db #(int)::set(null,"*","PORT_534_COUNT",port_count[534]);
       uvm_config_db #(int)::set(null,"*","PORT_535_COUNT",port_count[535]);
       uvm_config_db #(int)::set(null,"*","PORT_536_COUNT",port_count[536]);
       uvm_config_db #(int)::set(null,"*","PORT_537_COUNT",port_count[537]);
       uvm_config_db #(int)::set(null,"*","PORT_538_COUNT",port_count[538]);
       uvm_config_db #(int)::set(null,"*","PORT_539_COUNT",port_count[539]);
       uvm_config_db #(int)::set(null,"*","PORT_540_COUNT",port_count[540]);
       uvm_config_db #(int)::set(null,"*","PORT_541_COUNT",port_count[541]);
       uvm_config_db #(int)::set(null,"*","PORT_542_COUNT",port_count[542]);
       uvm_config_db #(int)::set(null,"*","PORT_543_COUNT",port_count[543]);
       uvm_config_db #(int)::set(null,"*","PORT_544_COUNT",port_count[544]);
       uvm_config_db #(int)::set(null,"*","PORT_545_COUNT",port_count[545]);
       uvm_config_db #(int)::set(null,"*","PORT_546_COUNT",port_count[546]);
       uvm_config_db #(int)::set(null,"*","PORT_547_COUNT",port_count[547]);
       uvm_config_db #(int)::set(null,"*","PORT_548_COUNT",port_count[548]);
       uvm_config_db #(int)::set(null,"*","PORT_549_COUNT",port_count[549]);
       uvm_config_db #(int)::set(null,"*","PORT_550_COUNT",port_count[550]);
       uvm_config_db #(int)::set(null,"*","PORT_551_COUNT",port_count[551]);
       uvm_config_db #(int)::set(null,"*","PORT_552_COUNT",port_count[552]);
       uvm_config_db #(int)::set(null,"*","PORT_553_COUNT",port_count[553]);
       uvm_config_db #(int)::set(null,"*","PORT_554_COUNT",port_count[554]);
       uvm_config_db #(int)::set(null,"*","PORT_555_COUNT",port_count[555]);
       uvm_config_db #(int)::set(null,"*","PORT_556_COUNT",port_count[556]);
       uvm_config_db #(int)::set(null,"*","PORT_557_COUNT",port_count[557]);
       uvm_config_db #(int)::set(null,"*","PORT_558_COUNT",port_count[558]);
       uvm_config_db #(int)::set(null,"*","PORT_559_COUNT",port_count[559]);
       uvm_config_db #(int)::set(null,"*","PORT_560_COUNT",port_count[560]);
       uvm_config_db #(int)::set(null,"*","PORT_561_COUNT",port_count[561]);
       uvm_config_db #(int)::set(null,"*","PORT_562_COUNT",port_count[562]);
       uvm_config_db #(int)::set(null,"*","PORT_563_COUNT",port_count[563]);
       uvm_config_db #(int)::set(null,"*","PORT_564_COUNT",port_count[564]);
       uvm_config_db #(int)::set(null,"*","PORT_565_COUNT",port_count[565]);
       uvm_config_db #(int)::set(null,"*","PORT_566_COUNT",port_count[566]);
       uvm_config_db #(int)::set(null,"*","PORT_567_COUNT",port_count[567]);
       uvm_config_db #(int)::set(null,"*","PORT_568_COUNT",port_count[568]);
       uvm_config_db #(int)::set(null,"*","PORT_569_COUNT",port_count[569]);
       uvm_config_db #(int)::set(null,"*","PORT_570_COUNT",port_count[570]);
       uvm_config_db #(int)::set(null,"*","PORT_571_COUNT",port_count[571]);
       uvm_config_db #(int)::set(null,"*","PORT_572_COUNT",port_count[572]);
       uvm_config_db #(int)::set(null,"*","PORT_573_COUNT",port_count[573]);
       uvm_config_db #(int)::set(null,"*","PORT_574_COUNT",port_count[574]);
       uvm_config_db #(int)::set(null,"*","PORT_575_COUNT",port_count[575]);
       uvm_config_db #(int)::set(null,"*","PORT_576_COUNT",port_count[576]);
       uvm_config_db #(int)::set(null,"*","PORT_577_COUNT",port_count[577]);
       uvm_config_db #(int)::set(null,"*","PORT_578_COUNT",port_count[578]);
       uvm_config_db #(int)::set(null,"*","PORT_579_COUNT",port_count[579]);
       uvm_config_db #(int)::set(null,"*","PORT_580_COUNT",port_count[580]);
       uvm_config_db #(int)::set(null,"*","PORT_581_COUNT",port_count[581]);
       uvm_config_db #(int)::set(null,"*","PORT_582_COUNT",port_count[582]);
       uvm_config_db #(int)::set(null,"*","PORT_583_COUNT",port_count[583]);
       uvm_config_db #(int)::set(null,"*","PORT_584_COUNT",port_count[584]);
       uvm_config_db #(int)::set(null,"*","PORT_585_COUNT",port_count[585]);
       uvm_config_db #(int)::set(null,"*","PORT_586_COUNT",port_count[586]);
       uvm_config_db #(int)::set(null,"*","PORT_587_COUNT",port_count[587]);
       uvm_config_db #(int)::set(null,"*","PORT_588_COUNT",port_count[588]);
       uvm_config_db #(int)::set(null,"*","PORT_589_COUNT",port_count[589]);
       uvm_config_db #(int)::set(null,"*","PORT_590_COUNT",port_count[590]);
       uvm_config_db #(int)::set(null,"*","PORT_591_COUNT",port_count[591]);
       uvm_config_db #(int)::set(null,"*","PORT_592_COUNT",port_count[592]);
       uvm_config_db #(int)::set(null,"*","PORT_593_COUNT",port_count[593]);
       uvm_config_db #(int)::set(null,"*","PORT_594_COUNT",port_count[594]);
       uvm_config_db #(int)::set(null,"*","PORT_595_COUNT",port_count[595]);
       uvm_config_db #(int)::set(null,"*","PORT_596_COUNT",port_count[596]);
       uvm_config_db #(int)::set(null,"*","PORT_597_COUNT",port_count[597]);
       uvm_config_db #(int)::set(null,"*","PORT_598_COUNT",port_count[598]);
       uvm_config_db #(int)::set(null,"*","PORT_599_COUNT",port_count[599]);
       uvm_config_db #(int)::set(null,"*","PORT_600_COUNT",port_count[600]);
       uvm_config_db #(int)::set(null,"*","PORT_601_COUNT",port_count[601]);
       uvm_config_db #(int)::set(null,"*","PORT_602_COUNT",port_count[602]);
       uvm_config_db #(int)::set(null,"*","PORT_603_COUNT",port_count[603]);
       uvm_config_db #(int)::set(null,"*","PORT_604_COUNT",port_count[604]);
       uvm_config_db #(int)::set(null,"*","PORT_605_COUNT",port_count[605]);
       uvm_config_db #(int)::set(null,"*","PORT_606_COUNT",port_count[606]);
       uvm_config_db #(int)::set(null,"*","PORT_607_COUNT",port_count[607]);
       uvm_config_db #(int)::set(null,"*","PORT_608_COUNT",port_count[608]);
       uvm_config_db #(int)::set(null,"*","PORT_609_COUNT",port_count[609]);
       uvm_config_db #(int)::set(null,"*","PORT_610_COUNT",port_count[610]);
       uvm_config_db #(int)::set(null,"*","PORT_611_COUNT",port_count[611]);
       uvm_config_db #(int)::set(null,"*","PORT_612_COUNT",port_count[612]);
       uvm_config_db #(int)::set(null,"*","PORT_613_COUNT",port_count[613]);
       uvm_config_db #(int)::set(null,"*","PORT_614_COUNT",port_count[614]);
       uvm_config_db #(int)::set(null,"*","PORT_615_COUNT",port_count[615]);
       uvm_config_db #(int)::set(null,"*","PORT_616_COUNT",port_count[616]);
       uvm_config_db #(int)::set(null,"*","PORT_617_COUNT",port_count[617]);
       uvm_config_db #(int)::set(null,"*","PORT_618_COUNT",port_count[618]);
       uvm_config_db #(int)::set(null,"*","PORT_619_COUNT",port_count[619]);
       uvm_config_db #(int)::set(null,"*","PORT_620_COUNT",port_count[620]);
       uvm_config_db #(int)::set(null,"*","PORT_621_COUNT",port_count[621]);
       uvm_config_db #(int)::set(null,"*","PORT_622_COUNT",port_count[622]);
       uvm_config_db #(int)::set(null,"*","PORT_623_COUNT",port_count[623]);
       uvm_config_db #(int)::set(null,"*","PORT_624_COUNT",port_count[624]);
       uvm_config_db #(int)::set(null,"*","PORT_625_COUNT",port_count[625]);
       uvm_config_db #(int)::set(null,"*","PORT_626_COUNT",port_count[626]);
       uvm_config_db #(int)::set(null,"*","PORT_627_COUNT",port_count[627]);
       uvm_config_db #(int)::set(null,"*","PORT_628_COUNT",port_count[628]);
       uvm_config_db #(int)::set(null,"*","PORT_629_COUNT",port_count[629]);
       uvm_config_db #(int)::set(null,"*","PORT_630_COUNT",port_count[630]);
       uvm_config_db #(int)::set(null,"*","PORT_631_COUNT",port_count[631]);
       uvm_config_db #(int)::set(null,"*","PORT_632_COUNT",port_count[632]);
       uvm_config_db #(int)::set(null,"*","PORT_633_COUNT",port_count[633]);
       uvm_config_db #(int)::set(null,"*","PORT_634_COUNT",port_count[634]);
       uvm_config_db #(int)::set(null,"*","PORT_635_COUNT",port_count[635]);
       uvm_config_db #(int)::set(null,"*","PORT_636_COUNT",port_count[636]);
       uvm_config_db #(int)::set(null,"*","PORT_637_COUNT",port_count[637]);
       uvm_config_db #(int)::set(null,"*","PORT_638_COUNT",port_count[638]);
       uvm_config_db #(int)::set(null,"*","PORT_639_COUNT",port_count[639]);
       uvm_config_db #(int)::set(null,"*","PORT_640_COUNT",port_count[640]);
       uvm_config_db #(int)::set(null,"*","PORT_641_COUNT",port_count[641]);
       uvm_config_db #(int)::set(null,"*","PORT_642_COUNT",port_count[642]);
       uvm_config_db #(int)::set(null,"*","PORT_643_COUNT",port_count[643]);
       uvm_config_db #(int)::set(null,"*","PORT_644_COUNT",port_count[644]);
       uvm_config_db #(int)::set(null,"*","PORT_645_COUNT",port_count[645]);
       uvm_config_db #(int)::set(null,"*","PORT_646_COUNT",port_count[646]);
       uvm_config_db #(int)::set(null,"*","PORT_647_COUNT",port_count[647]);
       uvm_config_db #(int)::set(null,"*","PORT_648_COUNT",port_count[648]);
       uvm_config_db #(int)::set(null,"*","PORT_649_COUNT",port_count[649]);
       uvm_config_db #(int)::set(null,"*","PORT_650_COUNT",port_count[650]);
       uvm_config_db #(int)::set(null,"*","PORT_651_COUNT",port_count[651]);
       uvm_config_db #(int)::set(null,"*","PORT_652_COUNT",port_count[652]);
       uvm_config_db #(int)::set(null,"*","PORT_653_COUNT",port_count[653]);
       uvm_config_db #(int)::set(null,"*","PORT_654_COUNT",port_count[654]);
       uvm_config_db #(int)::set(null,"*","PORT_655_COUNT",port_count[655]);
       uvm_config_db #(int)::set(null,"*","PORT_656_COUNT",port_count[656]);
       uvm_config_db #(int)::set(null,"*","PORT_657_COUNT",port_count[657]);
       uvm_config_db #(int)::set(null,"*","PORT_658_COUNT",port_count[658]);
       uvm_config_db #(int)::set(null,"*","PORT_659_COUNT",port_count[659]);
       uvm_config_db #(int)::set(null,"*","PORT_660_COUNT",port_count[660]);
       uvm_config_db #(int)::set(null,"*","PORT_661_COUNT",port_count[661]);
       uvm_config_db #(int)::set(null,"*","PORT_662_COUNT",port_count[662]);
       uvm_config_db #(int)::set(null,"*","PORT_663_COUNT",port_count[663]);
       uvm_config_db #(int)::set(null,"*","PORT_664_COUNT",port_count[664]);
       uvm_config_db #(int)::set(null,"*","PORT_665_COUNT",port_count[665]);
       uvm_config_db #(int)::set(null,"*","PORT_666_COUNT",port_count[666]);
       uvm_config_db #(int)::set(null,"*","PORT_667_COUNT",port_count[667]);
       uvm_config_db #(int)::set(null,"*","PORT_668_COUNT",port_count[668]);
       uvm_config_db #(int)::set(null,"*","PORT_669_COUNT",port_count[669]);
       uvm_config_db #(int)::set(null,"*","PORT_670_COUNT",port_count[670]);
       uvm_config_db #(int)::set(null,"*","PORT_671_COUNT",port_count[671]);
       uvm_config_db #(int)::set(null,"*","PORT_672_COUNT",port_count[672]);
       uvm_config_db #(int)::set(null,"*","PORT_673_COUNT",port_count[673]);
       uvm_config_db #(int)::set(null,"*","PORT_674_COUNT",port_count[674]);
       uvm_config_db #(int)::set(null,"*","PORT_675_COUNT",port_count[675]);
       uvm_config_db #(int)::set(null,"*","PORT_676_COUNT",port_count[676]);
       uvm_config_db #(int)::set(null,"*","PORT_677_COUNT",port_count[677]);
       uvm_config_db #(int)::set(null,"*","PORT_678_COUNT",port_count[678]);
       uvm_config_db #(int)::set(null,"*","PORT_679_COUNT",port_count[679]);
       uvm_config_db #(int)::set(null,"*","PORT_680_COUNT",port_count[680]);
       uvm_config_db #(int)::set(null,"*","PORT_681_COUNT",port_count[681]);
       uvm_config_db #(int)::set(null,"*","PORT_682_COUNT",port_count[682]);
       uvm_config_db #(int)::set(null,"*","PORT_683_COUNT",port_count[683]);
       uvm_config_db #(int)::set(null,"*","PORT_684_COUNT",port_count[684]);
       uvm_config_db #(int)::set(null,"*","PORT_685_COUNT",port_count[685]);
       uvm_config_db #(int)::set(null,"*","PORT_686_COUNT",port_count[686]);
       uvm_config_db #(int)::set(null,"*","PORT_687_COUNT",port_count[687]);
       uvm_config_db #(int)::set(null,"*","PORT_688_COUNT",port_count[688]);
       uvm_config_db #(int)::set(null,"*","PORT_689_COUNT",port_count[689]);
       uvm_config_db #(int)::set(null,"*","PORT_690_COUNT",port_count[690]);
       uvm_config_db #(int)::set(null,"*","PORT_691_COUNT",port_count[691]);
       uvm_config_db #(int)::set(null,"*","PORT_692_COUNT",port_count[692]);
       uvm_config_db #(int)::set(null,"*","PORT_693_COUNT",port_count[693]);
       uvm_config_db #(int)::set(null,"*","PORT_694_COUNT",port_count[694]);
       uvm_config_db #(int)::set(null,"*","PORT_695_COUNT",port_count[695]);
       uvm_config_db #(int)::set(null,"*","PORT_696_COUNT",port_count[696]);
       uvm_config_db #(int)::set(null,"*","PORT_697_COUNT",port_count[697]);
       uvm_config_db #(int)::set(null,"*","PORT_698_COUNT",port_count[698]);
       uvm_config_db #(int)::set(null,"*","PORT_699_COUNT",port_count[699]);
       uvm_config_db #(int)::set(null,"*","PORT_700_COUNT",port_count[700]);
       uvm_config_db #(int)::set(null,"*","PORT_701_COUNT",port_count[701]);
       uvm_config_db #(int)::set(null,"*","PORT_702_COUNT",port_count[702]);
       uvm_config_db #(int)::set(null,"*","PORT_703_COUNT",port_count[703]);
       uvm_config_db #(int)::set(null,"*","PORT_704_COUNT",port_count[704]);
       uvm_config_db #(int)::set(null,"*","PORT_705_COUNT",port_count[705]);
       uvm_config_db #(int)::set(null,"*","PORT_706_COUNT",port_count[706]);
       uvm_config_db #(int)::set(null,"*","PORT_707_COUNT",port_count[707]);
       uvm_config_db #(int)::set(null,"*","PORT_708_COUNT",port_count[708]);
       uvm_config_db #(int)::set(null,"*","PORT_709_COUNT",port_count[709]);
       uvm_config_db #(int)::set(null,"*","PORT_710_COUNT",port_count[710]);
       uvm_config_db #(int)::set(null,"*","PORT_711_COUNT",port_count[711]);
       uvm_config_db #(int)::set(null,"*","PORT_712_COUNT",port_count[712]);
       uvm_config_db #(int)::set(null,"*","PORT_713_COUNT",port_count[713]);
       uvm_config_db #(int)::set(null,"*","PORT_714_COUNT",port_count[714]);
       uvm_config_db #(int)::set(null,"*","PORT_715_COUNT",port_count[715]);
       uvm_config_db #(int)::set(null,"*","PORT_716_COUNT",port_count[716]);
       uvm_config_db #(int)::set(null,"*","PORT_717_COUNT",port_count[717]);
       uvm_config_db #(int)::set(null,"*","PORT_718_COUNT",port_count[718]);
       uvm_config_db #(int)::set(null,"*","PORT_719_COUNT",port_count[719]);
       uvm_config_db #(int)::set(null,"*","PORT_720_COUNT",port_count[720]);
       uvm_config_db #(int)::set(null,"*","PORT_721_COUNT",port_count[721]);
       uvm_config_db #(int)::set(null,"*","PORT_722_COUNT",port_count[722]);
       uvm_config_db #(int)::set(null,"*","PORT_723_COUNT",port_count[723]);
       uvm_config_db #(int)::set(null,"*","PORT_724_COUNT",port_count[724]);
       uvm_config_db #(int)::set(null,"*","PORT_725_COUNT",port_count[725]);
       uvm_config_db #(int)::set(null,"*","PORT_726_COUNT",port_count[726]);
       uvm_config_db #(int)::set(null,"*","PORT_727_COUNT",port_count[727]);
       uvm_config_db #(int)::set(null,"*","PORT_728_COUNT",port_count[728]);
       uvm_config_db #(int)::set(null,"*","PORT_729_COUNT",port_count[729]);
       uvm_config_db #(int)::set(null,"*","PORT_730_COUNT",port_count[730]);
       uvm_config_db #(int)::set(null,"*","PORT_731_COUNT",port_count[731]);
       uvm_config_db #(int)::set(null,"*","PORT_732_COUNT",port_count[732]);
       uvm_config_db #(int)::set(null,"*","PORT_733_COUNT",port_count[733]);
       uvm_config_db #(int)::set(null,"*","PORT_734_COUNT",port_count[734]);
       uvm_config_db #(int)::set(null,"*","PORT_735_COUNT",port_count[735]);
       uvm_config_db #(int)::set(null,"*","PORT_736_COUNT",port_count[736]);
       uvm_config_db #(int)::set(null,"*","PORT_737_COUNT",port_count[737]);
       uvm_config_db #(int)::set(null,"*","PORT_738_COUNT",port_count[738]);
       uvm_config_db #(int)::set(null,"*","PORT_739_COUNT",port_count[739]);
       uvm_config_db #(int)::set(null,"*","PORT_740_COUNT",port_count[740]);
       uvm_config_db #(int)::set(null,"*","PORT_741_COUNT",port_count[741]);
       uvm_config_db #(int)::set(null,"*","PORT_742_COUNT",port_count[742]);
       uvm_config_db #(int)::set(null,"*","PORT_743_COUNT",port_count[743]);
       uvm_config_db #(int)::set(null,"*","PORT_744_COUNT",port_count[744]);
       uvm_config_db #(int)::set(null,"*","PORT_745_COUNT",port_count[745]);
       uvm_config_db #(int)::set(null,"*","PORT_746_COUNT",port_count[746]);
       uvm_config_db #(int)::set(null,"*","PORT_747_COUNT",port_count[747]);
       uvm_config_db #(int)::set(null,"*","PORT_748_COUNT",port_count[748]);
       uvm_config_db #(int)::set(null,"*","PORT_749_COUNT",port_count[749]);
       uvm_config_db #(int)::set(null,"*","PORT_750_COUNT",port_count[750]);
       uvm_config_db #(int)::set(null,"*","PORT_751_COUNT",port_count[751]);
       uvm_config_db #(int)::set(null,"*","PORT_752_COUNT",port_count[752]);
       uvm_config_db #(int)::set(null,"*","PORT_753_COUNT",port_count[753]);
       uvm_config_db #(int)::set(null,"*","PORT_754_COUNT",port_count[754]);
       uvm_config_db #(int)::set(null,"*","PORT_755_COUNT",port_count[755]);
       uvm_config_db #(int)::set(null,"*","PORT_756_COUNT",port_count[756]);
       uvm_config_db #(int)::set(null,"*","PORT_757_COUNT",port_count[757]);
       uvm_config_db #(int)::set(null,"*","PORT_758_COUNT",port_count[758]);
       uvm_config_db #(int)::set(null,"*","PORT_759_COUNT",port_count[759]);
       uvm_config_db #(int)::set(null,"*","PORT_760_COUNT",port_count[760]);
       uvm_config_db #(int)::set(null,"*","PORT_761_COUNT",port_count[761]);
       uvm_config_db #(int)::set(null,"*","PORT_762_COUNT",port_count[762]);
       uvm_config_db #(int)::set(null,"*","PORT_763_COUNT",port_count[763]);
       uvm_config_db #(int)::set(null,"*","PORT_764_COUNT",port_count[764]);
       uvm_config_db #(int)::set(null,"*","PORT_765_COUNT",port_count[765]);
       uvm_config_db #(int)::set(null,"*","PORT_766_COUNT",port_count[766]);
       uvm_config_db #(int)::set(null,"*","PORT_767_COUNT",port_count[767]);
       uvm_config_db #(int)::set(null,"*","PORT_768_COUNT",port_count[768]);
       uvm_config_db #(int)::set(null,"*","PORT_769_COUNT",port_count[769]);
       uvm_config_db #(int)::set(null,"*","PORT_770_COUNT",port_count[770]);
       uvm_config_db #(int)::set(null,"*","PORT_771_COUNT",port_count[771]);
       uvm_config_db #(int)::set(null,"*","PORT_772_COUNT",port_count[772]);
       uvm_config_db #(int)::set(null,"*","PORT_773_COUNT",port_count[773]);
       uvm_config_db #(int)::set(null,"*","PORT_774_COUNT",port_count[774]);
       uvm_config_db #(int)::set(null,"*","PORT_775_COUNT",port_count[775]);
       uvm_config_db #(int)::set(null,"*","PORT_776_COUNT",port_count[776]);
       uvm_config_db #(int)::set(null,"*","PORT_777_COUNT",port_count[777]);
       uvm_config_db #(int)::set(null,"*","PORT_778_COUNT",port_count[778]);
       uvm_config_db #(int)::set(null,"*","PORT_779_COUNT",port_count[779]);
       uvm_config_db #(int)::set(null,"*","PORT_780_COUNT",port_count[780]);
       uvm_config_db #(int)::set(null,"*","PORT_781_COUNT",port_count[781]);
       uvm_config_db #(int)::set(null,"*","PORT_782_COUNT",port_count[782]);
       uvm_config_db #(int)::set(null,"*","PORT_783_COUNT",port_count[783]);
       uvm_config_db #(int)::set(null,"*","PORT_784_COUNT",port_count[784]);
       uvm_config_db #(int)::set(null,"*","PORT_785_COUNT",port_count[785]);
       uvm_config_db #(int)::set(null,"*","PORT_786_COUNT",port_count[786]);
       uvm_config_db #(int)::set(null,"*","PORT_787_COUNT",port_count[787]);
       uvm_config_db #(int)::set(null,"*","PORT_788_COUNT",port_count[788]);
       uvm_config_db #(int)::set(null,"*","PORT_789_COUNT",port_count[789]);
       uvm_config_db #(int)::set(null,"*","PORT_790_COUNT",port_count[790]);
       uvm_config_db #(int)::set(null,"*","PORT_791_COUNT",port_count[791]);
       uvm_config_db #(int)::set(null,"*","PORT_792_COUNT",port_count[792]);
       uvm_config_db #(int)::set(null,"*","PORT_793_COUNT",port_count[793]);
       uvm_config_db #(int)::set(null,"*","PORT_794_COUNT",port_count[794]);
       uvm_config_db #(int)::set(null,"*","PORT_795_COUNT",port_count[795]);
       uvm_config_db #(int)::set(null,"*","PORT_796_COUNT",port_count[796]);
       uvm_config_db #(int)::set(null,"*","PORT_797_COUNT",port_count[797]);
       uvm_config_db #(int)::set(null,"*","PORT_798_COUNT",port_count[798]);
       uvm_config_db #(int)::set(null,"*","PORT_799_COUNT",port_count[799]);
       uvm_config_db #(int)::set(null,"*","PORT_800_COUNT",port_count[800]);
       uvm_config_db #(int)::set(null,"*","PORT_801_COUNT",port_count[801]);
       uvm_config_db #(int)::set(null,"*","PORT_802_COUNT",port_count[802]);
       uvm_config_db #(int)::set(null,"*","PORT_803_COUNT",port_count[803]);
       uvm_config_db #(int)::set(null,"*","PORT_804_COUNT",port_count[804]);
       uvm_config_db #(int)::set(null,"*","PORT_805_COUNT",port_count[805]);
       uvm_config_db #(int)::set(null,"*","PORT_806_COUNT",port_count[806]);
       uvm_config_db #(int)::set(null,"*","PORT_807_COUNT",port_count[807]);
       uvm_config_db #(int)::set(null,"*","PORT_808_COUNT",port_count[808]);
       uvm_config_db #(int)::set(null,"*","PORT_809_COUNT",port_count[809]);
       uvm_config_db #(int)::set(null,"*","PORT_810_COUNT",port_count[810]);
       uvm_config_db #(int)::set(null,"*","PORT_811_COUNT",port_count[811]);
       uvm_config_db #(int)::set(null,"*","PORT_812_COUNT",port_count[812]);
       uvm_config_db #(int)::set(null,"*","PORT_813_COUNT",port_count[813]);
       uvm_config_db #(int)::set(null,"*","PORT_814_COUNT",port_count[814]);
       uvm_config_db #(int)::set(null,"*","PORT_815_COUNT",port_count[815]);
       uvm_config_db #(int)::set(null,"*","PORT_816_COUNT",port_count[816]);
       uvm_config_db #(int)::set(null,"*","PORT_817_COUNT",port_count[817]);
       uvm_config_db #(int)::set(null,"*","PORT_818_COUNT",port_count[818]);
       uvm_config_db #(int)::set(null,"*","PORT_819_COUNT",port_count[819]);
       uvm_config_db #(int)::set(null,"*","PORT_820_COUNT",port_count[820]);
       uvm_config_db #(int)::set(null,"*","PORT_821_COUNT",port_count[821]);
       uvm_config_db #(int)::set(null,"*","PORT_822_COUNT",port_count[822]);
       uvm_config_db #(int)::set(null,"*","PORT_823_COUNT",port_count[823]);
       uvm_config_db #(int)::set(null,"*","PORT_824_COUNT",port_count[824]);
       uvm_config_db #(int)::set(null,"*","PORT_825_COUNT",port_count[825]);
       uvm_config_db #(int)::set(null,"*","PORT_826_COUNT",port_count[826]);
       uvm_config_db #(int)::set(null,"*","PORT_827_COUNT",port_count[827]);
       uvm_config_db #(int)::set(null,"*","PORT_828_COUNT",port_count[828]);
       uvm_config_db #(int)::set(null,"*","PORT_829_COUNT",port_count[829]);
       uvm_config_db #(int)::set(null,"*","PORT_830_COUNT",port_count[830]);
       uvm_config_db #(int)::set(null,"*","PORT_831_COUNT",port_count[831]);
       uvm_config_db #(int)::set(null,"*","PORT_832_COUNT",port_count[832]);
       uvm_config_db #(int)::set(null,"*","PORT_833_COUNT",port_count[833]);
       uvm_config_db #(int)::set(null,"*","PORT_834_COUNT",port_count[834]);
       uvm_config_db #(int)::set(null,"*","PORT_835_COUNT",port_count[835]);
       uvm_config_db #(int)::set(null,"*","PORT_836_COUNT",port_count[836]);
       uvm_config_db #(int)::set(null,"*","PORT_837_COUNT",port_count[837]);
       uvm_config_db #(int)::set(null,"*","PORT_838_COUNT",port_count[838]);
       uvm_config_db #(int)::set(null,"*","PORT_839_COUNT",port_count[839]);
       uvm_config_db #(int)::set(null,"*","PORT_840_COUNT",port_count[840]);
       uvm_config_db #(int)::set(null,"*","PORT_841_COUNT",port_count[841]);
       uvm_config_db #(int)::set(null,"*","PORT_842_COUNT",port_count[842]);
       uvm_config_db #(int)::set(null,"*","PORT_843_COUNT",port_count[843]);
       uvm_config_db #(int)::set(null,"*","PORT_844_COUNT",port_count[844]);
       uvm_config_db #(int)::set(null,"*","PORT_845_COUNT",port_count[845]);
       uvm_config_db #(int)::set(null,"*","PORT_846_COUNT",port_count[846]);
       uvm_config_db #(int)::set(null,"*","PORT_847_COUNT",port_count[847]);
       uvm_config_db #(int)::set(null,"*","PORT_848_COUNT",port_count[848]);
       uvm_config_db #(int)::set(null,"*","PORT_849_COUNT",port_count[849]);
       uvm_config_db #(int)::set(null,"*","PORT_850_COUNT",port_count[850]);
       uvm_config_db #(int)::set(null,"*","PORT_851_COUNT",port_count[851]);
       uvm_config_db #(int)::set(null,"*","PORT_852_COUNT",port_count[852]);
       uvm_config_db #(int)::set(null,"*","PORT_853_COUNT",port_count[853]);
       uvm_config_db #(int)::set(null,"*","PORT_854_COUNT",port_count[854]);
       uvm_config_db #(int)::set(null,"*","PORT_855_COUNT",port_count[855]);
       uvm_config_db #(int)::set(null,"*","PORT_856_COUNT",port_count[856]);
       uvm_config_db #(int)::set(null,"*","PORT_857_COUNT",port_count[857]);
       uvm_config_db #(int)::set(null,"*","PORT_858_COUNT",port_count[858]);
       uvm_config_db #(int)::set(null,"*","PORT_859_COUNT",port_count[859]);
       uvm_config_db #(int)::set(null,"*","PORT_860_COUNT",port_count[860]);
       uvm_config_db #(int)::set(null,"*","PORT_861_COUNT",port_count[861]);
       uvm_config_db #(int)::set(null,"*","PORT_862_COUNT",port_count[862]);
       uvm_config_db #(int)::set(null,"*","PORT_863_COUNT",port_count[863]);
       uvm_config_db #(int)::set(null,"*","PORT_864_COUNT",port_count[864]);
       uvm_config_db #(int)::set(null,"*","PORT_865_COUNT",port_count[865]);
       uvm_config_db #(int)::set(null,"*","PORT_866_COUNT",port_count[866]);
       uvm_config_db #(int)::set(null,"*","PORT_867_COUNT",port_count[867]);
       uvm_config_db #(int)::set(null,"*","PORT_868_COUNT",port_count[868]);
       uvm_config_db #(int)::set(null,"*","PORT_869_COUNT",port_count[869]);
       uvm_config_db #(int)::set(null,"*","PORT_870_COUNT",port_count[870]);
       uvm_config_db #(int)::set(null,"*","PORT_871_COUNT",port_count[871]);
       uvm_config_db #(int)::set(null,"*","PORT_872_COUNT",port_count[872]);
       uvm_config_db #(int)::set(null,"*","PORT_873_COUNT",port_count[873]);
       uvm_config_db #(int)::set(null,"*","PORT_874_COUNT",port_count[874]);
       uvm_config_db #(int)::set(null,"*","PORT_875_COUNT",port_count[875]);
       uvm_config_db #(int)::set(null,"*","PORT_876_COUNT",port_count[876]);
       uvm_config_db #(int)::set(null,"*","PORT_877_COUNT",port_count[877]);
       uvm_config_db #(int)::set(null,"*","PORT_878_COUNT",port_count[878]);
       uvm_config_db #(int)::set(null,"*","PORT_879_COUNT",port_count[879]);
       uvm_config_db #(int)::set(null,"*","PORT_880_COUNT",port_count[880]);
       uvm_config_db #(int)::set(null,"*","PORT_881_COUNT",port_count[881]);
       uvm_config_db #(int)::set(null,"*","PORT_882_COUNT",port_count[882]);
       uvm_config_db #(int)::set(null,"*","PORT_883_COUNT",port_count[883]);
       uvm_config_db #(int)::set(null,"*","PORT_884_COUNT",port_count[884]);
       uvm_config_db #(int)::set(null,"*","PORT_885_COUNT",port_count[885]);
       uvm_config_db #(int)::set(null,"*","PORT_886_COUNT",port_count[886]);
       uvm_config_db #(int)::set(null,"*","PORT_887_COUNT",port_count[887]);
       uvm_config_db #(int)::set(null,"*","PORT_888_COUNT",port_count[888]);
       uvm_config_db #(int)::set(null,"*","PORT_889_COUNT",port_count[889]);
       uvm_config_db #(int)::set(null,"*","PORT_890_COUNT",port_count[890]);
       uvm_config_db #(int)::set(null,"*","PORT_891_COUNT",port_count[891]);
       uvm_config_db #(int)::set(null,"*","PORT_892_COUNT",port_count[892]);
       uvm_config_db #(int)::set(null,"*","PORT_893_COUNT",port_count[893]);
       uvm_config_db #(int)::set(null,"*","PORT_894_COUNT",port_count[894]);
       uvm_config_db #(int)::set(null,"*","PORT_895_COUNT",port_count[895]);
       uvm_config_db #(int)::set(null,"*","PORT_896_COUNT",port_count[896]);
       uvm_config_db #(int)::set(null,"*","PORT_897_COUNT",port_count[897]);
       uvm_config_db #(int)::set(null,"*","PORT_898_COUNT",port_count[898]);
       uvm_config_db #(int)::set(null,"*","PORT_899_COUNT",port_count[899]);
       uvm_config_db #(int)::set(null,"*","PORT_900_COUNT",port_count[900]);
       uvm_config_db #(int)::set(null,"*","PORT_901_COUNT",port_count[901]);
       uvm_config_db #(int)::set(null,"*","PORT_902_COUNT",port_count[902]);
       uvm_config_db #(int)::set(null,"*","PORT_903_COUNT",port_count[903]);
       uvm_config_db #(int)::set(null,"*","PORT_904_COUNT",port_count[904]);
       uvm_config_db #(int)::set(null,"*","PORT_905_COUNT",port_count[905]);
       uvm_config_db #(int)::set(null,"*","PORT_906_COUNT",port_count[906]);
       uvm_config_db #(int)::set(null,"*","PORT_907_COUNT",port_count[907]);
       uvm_config_db #(int)::set(null,"*","PORT_908_COUNT",port_count[908]);
       uvm_config_db #(int)::set(null,"*","PORT_909_COUNT",port_count[909]);
       uvm_config_db #(int)::set(null,"*","PORT_910_COUNT",port_count[910]);
       uvm_config_db #(int)::set(null,"*","PORT_911_COUNT",port_count[911]);
       uvm_config_db #(int)::set(null,"*","PORT_912_COUNT",port_count[912]);
       uvm_config_db #(int)::set(null,"*","PORT_913_COUNT",port_count[913]);
       uvm_config_db #(int)::set(null,"*","PORT_914_COUNT",port_count[914]);
       uvm_config_db #(int)::set(null,"*","PORT_915_COUNT",port_count[915]);
       uvm_config_db #(int)::set(null,"*","PORT_916_COUNT",port_count[916]);
       uvm_config_db #(int)::set(null,"*","PORT_917_COUNT",port_count[917]);
       uvm_config_db #(int)::set(null,"*","PORT_918_COUNT",port_count[918]);
       uvm_config_db #(int)::set(null,"*","PORT_919_COUNT",port_count[919]);
       uvm_config_db #(int)::set(null,"*","PORT_920_COUNT",port_count[920]);
       uvm_config_db #(int)::set(null,"*","PORT_921_COUNT",port_count[921]);
       uvm_config_db #(int)::set(null,"*","PORT_922_COUNT",port_count[922]);
       uvm_config_db #(int)::set(null,"*","PORT_923_COUNT",port_count[923]);
       uvm_config_db #(int)::set(null,"*","PORT_924_COUNT",port_count[924]);
       uvm_config_db #(int)::set(null,"*","PORT_925_COUNT",port_count[925]);
       uvm_config_db #(int)::set(null,"*","PORT_926_COUNT",port_count[926]);
       uvm_config_db #(int)::set(null,"*","PORT_927_COUNT",port_count[927]);
       uvm_config_db #(int)::set(null,"*","PORT_928_COUNT",port_count[928]);
       uvm_config_db #(int)::set(null,"*","PORT_929_COUNT",port_count[929]);
       uvm_config_db #(int)::set(null,"*","PORT_930_COUNT",port_count[930]);
       uvm_config_db #(int)::set(null,"*","PORT_931_COUNT",port_count[931]);
       uvm_config_db #(int)::set(null,"*","PORT_932_COUNT",port_count[932]);
       uvm_config_db #(int)::set(null,"*","PORT_933_COUNT",port_count[933]);
       uvm_config_db #(int)::set(null,"*","PORT_934_COUNT",port_count[934]);
       uvm_config_db #(int)::set(null,"*","PORT_935_COUNT",port_count[935]);
       uvm_config_db #(int)::set(null,"*","PORT_936_COUNT",port_count[936]);
       uvm_config_db #(int)::set(null,"*","PORT_937_COUNT",port_count[937]);
       uvm_config_db #(int)::set(null,"*","PORT_938_COUNT",port_count[938]);
       uvm_config_db #(int)::set(null,"*","PORT_939_COUNT",port_count[939]);
       uvm_config_db #(int)::set(null,"*","PORT_940_COUNT",port_count[940]);
       uvm_config_db #(int)::set(null,"*","PORT_941_COUNT",port_count[941]);
       uvm_config_db #(int)::set(null,"*","PORT_942_COUNT",port_count[942]);
       uvm_config_db #(int)::set(null,"*","PORT_943_COUNT",port_count[943]);
       uvm_config_db #(int)::set(null,"*","PORT_944_COUNT",port_count[944]);
       uvm_config_db #(int)::set(null,"*","PORT_945_COUNT",port_count[945]);
       uvm_config_db #(int)::set(null,"*","PORT_946_COUNT",port_count[946]);
       uvm_config_db #(int)::set(null,"*","PORT_947_COUNT",port_count[947]);
       uvm_config_db #(int)::set(null,"*","PORT_948_COUNT",port_count[948]);
       uvm_config_db #(int)::set(null,"*","PORT_949_COUNT",port_count[949]);
       uvm_config_db #(int)::set(null,"*","PORT_950_COUNT",port_count[950]);
       uvm_config_db #(int)::set(null,"*","PORT_951_COUNT",port_count[951]);
       uvm_config_db #(int)::set(null,"*","PORT_952_COUNT",port_count[952]);
       uvm_config_db #(int)::set(null,"*","PORT_953_COUNT",port_count[953]);
       uvm_config_db #(int)::set(null,"*","PORT_954_COUNT",port_count[954]);
       uvm_config_db #(int)::set(null,"*","PORT_955_COUNT",port_count[955]);
       uvm_config_db #(int)::set(null,"*","PORT_956_COUNT",port_count[956]);
       uvm_config_db #(int)::set(null,"*","PORT_957_COUNT",port_count[957]);
       uvm_config_db #(int)::set(null,"*","PORT_958_COUNT",port_count[958]);
       uvm_config_db #(int)::set(null,"*","PORT_959_COUNT",port_count[959]);
       uvm_config_db #(int)::set(null,"*","PORT_960_COUNT",port_count[960]);
       uvm_config_db #(int)::set(null,"*","PORT_961_COUNT",port_count[961]);
       uvm_config_db #(int)::set(null,"*","PORT_962_COUNT",port_count[962]);
       uvm_config_db #(int)::set(null,"*","PORT_963_COUNT",port_count[963]);
       uvm_config_db #(int)::set(null,"*","PORT_964_COUNT",port_count[964]);
       uvm_config_db #(int)::set(null,"*","PORT_965_COUNT",port_count[965]);
       uvm_config_db #(int)::set(null,"*","PORT_966_COUNT",port_count[966]);
       uvm_config_db #(int)::set(null,"*","PORT_967_COUNT",port_count[967]);
       uvm_config_db #(int)::set(null,"*","PORT_968_COUNT",port_count[968]);
       uvm_config_db #(int)::set(null,"*","PORT_969_COUNT",port_count[969]);
       uvm_config_db #(int)::set(null,"*","PORT_970_COUNT",port_count[970]);
       uvm_config_db #(int)::set(null,"*","PORT_971_COUNT",port_count[971]);
       uvm_config_db #(int)::set(null,"*","PORT_972_COUNT",port_count[972]);
       uvm_config_db #(int)::set(null,"*","PORT_973_COUNT",port_count[973]);
       uvm_config_db #(int)::set(null,"*","PORT_974_COUNT",port_count[974]);
       uvm_config_db #(int)::set(null,"*","PORT_975_COUNT",port_count[975]);
       uvm_config_db #(int)::set(null,"*","PORT_976_COUNT",port_count[976]);
       uvm_config_db #(int)::set(null,"*","PORT_977_COUNT",port_count[977]);
       uvm_config_db #(int)::set(null,"*","PORT_978_COUNT",port_count[978]);
       uvm_config_db #(int)::set(null,"*","PORT_979_COUNT",port_count[979]);
       uvm_config_db #(int)::set(null,"*","PORT_980_COUNT",port_count[980]);
       uvm_config_db #(int)::set(null,"*","PORT_981_COUNT",port_count[981]);
       uvm_config_db #(int)::set(null,"*","PORT_982_COUNT",port_count[982]);
       uvm_config_db #(int)::set(null,"*","PORT_983_COUNT",port_count[983]);
       uvm_config_db #(int)::set(null,"*","PORT_984_COUNT",port_count[984]);
       uvm_config_db #(int)::set(null,"*","PORT_985_COUNT",port_count[985]);
       uvm_config_db #(int)::set(null,"*","PORT_986_COUNT",port_count[986]);
       uvm_config_db #(int)::set(null,"*","PORT_987_COUNT",port_count[987]);
       uvm_config_db #(int)::set(null,"*","PORT_988_COUNT",port_count[988]);
       uvm_config_db #(int)::set(null,"*","PORT_989_COUNT",port_count[989]);
       uvm_config_db #(int)::set(null,"*","PORT_990_COUNT",port_count[990]);
       uvm_config_db #(int)::set(null,"*","PORT_991_COUNT",port_count[991]);
       uvm_config_db #(int)::set(null,"*","PORT_992_COUNT",port_count[992]);
       uvm_config_db #(int)::set(null,"*","PORT_993_COUNT",port_count[993]);
       uvm_config_db #(int)::set(null,"*","PORT_994_COUNT",port_count[994]);
       uvm_config_db #(int)::set(null,"*","PORT_995_COUNT",port_count[995]);
       uvm_config_db #(int)::set(null,"*","PORT_996_COUNT",port_count[996]);
       uvm_config_db #(int)::set(null,"*","PORT_997_COUNT",port_count[997]);
       uvm_config_db #(int)::set(null,"*","PORT_998_COUNT",port_count[998]);
       uvm_config_db #(int)::set(null,"*","PORT_999_COUNT",port_count[999]);
       uvm_config_db #(int)::set(null,"*","PORT_1000_COUNT",port_count[1000]);
       uvm_config_db #(int)::set(null,"*","PORT_1001_COUNT",port_count[1001]);
       uvm_config_db #(int)::set(null,"*","PORT_1002_COUNT",port_count[1002]);
       uvm_config_db #(int)::set(null,"*","PORT_1003_COUNT",port_count[1003]);
       uvm_config_db #(int)::set(null,"*","PORT_1004_COUNT",port_count[1004]);
       uvm_config_db #(int)::set(null,"*","PORT_1005_COUNT",port_count[1005]);
       uvm_config_db #(int)::set(null,"*","PORT_1006_COUNT",port_count[1006]);
       uvm_config_db #(int)::set(null,"*","PORT_1007_COUNT",port_count[1007]);
       uvm_config_db #(int)::set(null,"*","PORT_1008_COUNT",port_count[1008]);
       uvm_config_db #(int)::set(null,"*","PORT_1009_COUNT",port_count[1009]);
       uvm_config_db #(int)::set(null,"*","PORT_1010_COUNT",port_count[1010]);
       uvm_config_db #(int)::set(null,"*","PORT_1011_COUNT",port_count[1011]);
       uvm_config_db #(int)::set(null,"*","PORT_1012_COUNT",port_count[1012]);
       uvm_config_db #(int)::set(null,"*","PORT_1013_COUNT",port_count[1013]);
       uvm_config_db #(int)::set(null,"*","PORT_1014_COUNT",port_count[1014]);
       uvm_config_db #(int)::set(null,"*","PORT_1015_COUNT",port_count[1015]);
       uvm_config_db #(int)::set(null,"*","PORT_1016_COUNT",port_count[1016]);
       uvm_config_db #(int)::set(null,"*","PORT_1017_COUNT",port_count[1017]);
       uvm_config_db #(int)::set(null,"*","PORT_1018_COUNT",port_count[1018]);
       uvm_config_db #(int)::set(null,"*","PORT_1019_COUNT",port_count[1019]);
       uvm_config_db #(int)::set(null,"*","PORT_1020_COUNT",port_count[1020]);
       uvm_config_db #(int)::set(null,"*","PORT_1021_COUNT",port_count[1021]);
       uvm_config_db #(int)::set(null,"*","PORT_1022_COUNT",port_count[1022]);
       uvm_config_db #(int)::set(null,"*","PORT_1023_COUNT",port_count[1023]);
       uvm_config_db #(int)::set(null,"*","PORT_1024_COUNT",port_count[1024]);
       uvm_config_db #(int)::set(null,"*","PORT_1025_COUNT",port_count[1025]);
       uvm_config_db #(int)::set(null,"*","PORT_1026_COUNT",port_count[1026]);
       uvm_config_db #(int)::set(null,"*","PORT_1027_COUNT",port_count[1027]);
       uvm_config_db #(int)::set(null,"*","PORT_1028_COUNT",port_count[1028]);
       uvm_config_db #(int)::set(null,"*","PORT_1029_COUNT",port_count[1029]);
       uvm_config_db #(int)::set(null,"*","PORT_1030_COUNT",port_count[1030]);
       uvm_config_db #(int)::set(null,"*","PORT_1031_COUNT",port_count[1031]);
       uvm_config_db #(int)::set(null,"*","PORT_1032_COUNT",port_count[1032]);
       uvm_config_db #(int)::set(null,"*","PORT_1033_COUNT",port_count[1033]);
       uvm_config_db #(int)::set(null,"*","PORT_1034_COUNT",port_count[1034]);
       uvm_config_db #(int)::set(null,"*","PORT_1035_COUNT",port_count[1035]);
       uvm_config_db #(int)::set(null,"*","PORT_1036_COUNT",port_count[1036]);
       uvm_config_db #(int)::set(null,"*","PORT_1037_COUNT",port_count[1037]);
       uvm_config_db #(int)::set(null,"*","PORT_1038_COUNT",port_count[1038]);
       uvm_config_db #(int)::set(null,"*","PORT_1039_COUNT",port_count[1039]);
       uvm_config_db #(int)::set(null,"*","PORT_1040_COUNT",port_count[1040]);
       uvm_config_db #(int)::set(null,"*","PORT_1041_COUNT",port_count[1041]);
       uvm_config_db #(int)::set(null,"*","PORT_1042_COUNT",port_count[1042]);
       uvm_config_db #(int)::set(null,"*","PORT_1043_COUNT",port_count[1043]);
       uvm_config_db #(int)::set(null,"*","PORT_1044_COUNT",port_count[1044]);
       uvm_config_db #(int)::set(null,"*","PORT_1045_COUNT",port_count[1045]);
       uvm_config_db #(int)::set(null,"*","PORT_1046_COUNT",port_count[1046]);
       uvm_config_db #(int)::set(null,"*","PORT_1047_COUNT",port_count[1047]);
       uvm_config_db #(int)::set(null,"*","PORT_1048_COUNT",port_count[1048]);
       uvm_config_db #(int)::set(null,"*","PORT_1049_COUNT",port_count[1049]);
       uvm_config_db #(int)::set(null,"*","PORT_1050_COUNT",port_count[1050]);
       uvm_config_db #(int)::set(null,"*","PORT_1051_COUNT",port_count[1051]);
       uvm_config_db #(int)::set(null,"*","PORT_1052_COUNT",port_count[1052]);
       uvm_config_db #(int)::set(null,"*","PORT_1053_COUNT",port_count[1053]);
       uvm_config_db #(int)::set(null,"*","PORT_1054_COUNT",port_count[1054]);
       uvm_config_db #(int)::set(null,"*","PORT_1055_COUNT",port_count[1055]);
       uvm_config_db #(int)::set(null,"*","PORT_1056_COUNT",port_count[1056]);
       uvm_config_db #(int)::set(null,"*","PORT_1057_COUNT",port_count[1057]);
       uvm_config_db #(int)::set(null,"*","PORT_1058_COUNT",port_count[1058]);
       uvm_config_db #(int)::set(null,"*","PORT_1059_COUNT",port_count[1059]);
       uvm_config_db #(int)::set(null,"*","PORT_1060_COUNT",port_count[1060]);
       uvm_config_db #(int)::set(null,"*","PORT_1061_COUNT",port_count[1061]);
       uvm_config_db #(int)::set(null,"*","PORT_1062_COUNT",port_count[1062]);
       uvm_config_db #(int)::set(null,"*","PORT_1063_COUNT",port_count[1063]);
       uvm_config_db #(int)::set(null,"*","PORT_1064_COUNT",port_count[1064]);
       uvm_config_db #(int)::set(null,"*","PORT_1065_COUNT",port_count[1065]);
       uvm_config_db #(int)::set(null,"*","PORT_1066_COUNT",port_count[1066]);
       uvm_config_db #(int)::set(null,"*","PORT_1067_COUNT",port_count[1067]);
       uvm_config_db #(int)::set(null,"*","PORT_1068_COUNT",port_count[1068]);
       uvm_config_db #(int)::set(null,"*","PORT_1069_COUNT",port_count[1069]);
       uvm_config_db #(int)::set(null,"*","PORT_1070_COUNT",port_count[1070]);
       uvm_config_db #(int)::set(null,"*","PORT_1071_COUNT",port_count[1071]);
       uvm_config_db #(int)::set(null,"*","PORT_1072_COUNT",port_count[1072]);
       uvm_config_db #(int)::set(null,"*","PORT_1073_COUNT",port_count[1073]);
       uvm_config_db #(int)::set(null,"*","PORT_1074_COUNT",port_count[1074]);
       uvm_config_db #(int)::set(null,"*","PORT_1075_COUNT",port_count[1075]);
       uvm_config_db #(int)::set(null,"*","PORT_1076_COUNT",port_count[1076]);
       uvm_config_db #(int)::set(null,"*","PORT_1077_COUNT",port_count[1077]);
       uvm_config_db #(int)::set(null,"*","PORT_1078_COUNT",port_count[1078]);
       uvm_config_db #(int)::set(null,"*","PORT_1079_COUNT",port_count[1079]);
       uvm_config_db #(int)::set(null,"*","PORT_1080_COUNT",port_count[1080]);
       uvm_config_db #(int)::set(null,"*","PORT_1081_COUNT",port_count[1081]);
       uvm_config_db #(int)::set(null,"*","PORT_1082_COUNT",port_count[1082]);
       uvm_config_db #(int)::set(null,"*","PORT_1083_COUNT",port_count[1083]);
       uvm_config_db #(int)::set(null,"*","PORT_1084_COUNT",port_count[1084]);
       uvm_config_db #(int)::set(null,"*","PORT_1085_COUNT",port_count[1085]);
       uvm_config_db #(int)::set(null,"*","PORT_1086_COUNT",port_count[1086]);
       uvm_config_db #(int)::set(null,"*","PORT_1087_COUNT",port_count[1087]);
       uvm_config_db #(int)::set(null,"*","PORT_1088_COUNT",port_count[1088]);
       uvm_config_db #(int)::set(null,"*","PORT_1089_COUNT",port_count[1089]);
       uvm_config_db #(int)::set(null,"*","PORT_1090_COUNT",port_count[1090]);
       uvm_config_db #(int)::set(null,"*","PORT_1091_COUNT",port_count[1091]);
       uvm_config_db #(int)::set(null,"*","PORT_1092_COUNT",port_count[1092]);
       uvm_config_db #(int)::set(null,"*","PORT_1093_COUNT",port_count[1093]);
       uvm_config_db #(int)::set(null,"*","PORT_1094_COUNT",port_count[1094]);
       uvm_config_db #(int)::set(null,"*","PORT_1095_COUNT",port_count[1095]);
       uvm_config_db #(int)::set(null,"*","PORT_1096_COUNT",port_count[1096]);
       uvm_config_db #(int)::set(null,"*","PORT_1097_COUNT",port_count[1097]);
       uvm_config_db #(int)::set(null,"*","PORT_1098_COUNT",port_count[1098]);
       uvm_config_db #(int)::set(null,"*","PORT_1099_COUNT",port_count[1099]);
       uvm_config_db #(int)::set(null,"*","PORT_1100_COUNT",port_count[1100]);
       uvm_config_db #(int)::set(null,"*","PORT_1101_COUNT",port_count[1101]);
       uvm_config_db #(int)::set(null,"*","PORT_1102_COUNT",port_count[1102]);
       uvm_config_db #(int)::set(null,"*","PORT_1103_COUNT",port_count[1103]);
       uvm_config_db #(int)::set(null,"*","PORT_1104_COUNT",port_count[1104]);
       uvm_config_db #(int)::set(null,"*","PORT_1105_COUNT",port_count[1105]);
       uvm_config_db #(int)::set(null,"*","PORT_1106_COUNT",port_count[1106]);
       uvm_config_db #(int)::set(null,"*","PORT_1107_COUNT",port_count[1107]);
       uvm_config_db #(int)::set(null,"*","PORT_1108_COUNT",port_count[1108]);
       uvm_config_db #(int)::set(null,"*","PORT_1109_COUNT",port_count[1109]);
       uvm_config_db #(int)::set(null,"*","PORT_1110_COUNT",port_count[1110]);
       uvm_config_db #(int)::set(null,"*","PORT_1111_COUNT",port_count[1111]);
       uvm_config_db #(int)::set(null,"*","PORT_1112_COUNT",port_count[1112]);
       uvm_config_db #(int)::set(null,"*","PORT_1113_COUNT",port_count[1113]);
       uvm_config_db #(int)::set(null,"*","PORT_1114_COUNT",port_count[1114]);
       uvm_config_db #(int)::set(null,"*","PORT_1115_COUNT",port_count[1115]);
       uvm_config_db #(int)::set(null,"*","PORT_1116_COUNT",port_count[1116]);
       uvm_config_db #(int)::set(null,"*","PORT_1117_COUNT",port_count[1117]);
       uvm_config_db #(int)::set(null,"*","PORT_1118_COUNT",port_count[1118]);
       uvm_config_db #(int)::set(null,"*","PORT_1119_COUNT",port_count[1119]);
       uvm_config_db #(int)::set(null,"*","PORT_1120_COUNT",port_count[1120]);
       uvm_config_db #(int)::set(null,"*","PORT_1121_COUNT",port_count[1121]);
       uvm_config_db #(int)::set(null,"*","PORT_1122_COUNT",port_count[1122]);
       uvm_config_db #(int)::set(null,"*","PORT_1123_COUNT",port_count[1123]);
       uvm_config_db #(int)::set(null,"*","PORT_1124_COUNT",port_count[1124]);
       uvm_config_db #(int)::set(null,"*","PORT_1125_COUNT",port_count[1125]);
       uvm_config_db #(int)::set(null,"*","PORT_1126_COUNT",port_count[1126]);
       uvm_config_db #(int)::set(null,"*","PORT_1127_COUNT",port_count[1127]);
       uvm_config_db #(int)::set(null,"*","PORT_1128_COUNT",port_count[1128]);
       uvm_config_db #(int)::set(null,"*","PORT_1129_COUNT",port_count[1129]);
       uvm_config_db #(int)::set(null,"*","PORT_1130_COUNT",port_count[1130]);
       uvm_config_db #(int)::set(null,"*","PORT_1131_COUNT",port_count[1131]);
       uvm_config_db #(int)::set(null,"*","PORT_1132_COUNT",port_count[1132]);
       uvm_config_db #(int)::set(null,"*","PORT_1133_COUNT",port_count[1133]);
       uvm_config_db #(int)::set(null,"*","PORT_1134_COUNT",port_count[1134]);
       uvm_config_db #(int)::set(null,"*","PORT_1135_COUNT",port_count[1135]);
       uvm_config_db #(int)::set(null,"*","PORT_1136_COUNT",port_count[1136]);
       uvm_config_db #(int)::set(null,"*","PORT_1137_COUNT",port_count[1137]);
       uvm_config_db #(int)::set(null,"*","PORT_1138_COUNT",port_count[1138]);
       uvm_config_db #(int)::set(null,"*","PORT_1139_COUNT",port_count[1139]);
       uvm_config_db #(int)::set(null,"*","PORT_1140_COUNT",port_count[1140]);
       uvm_config_db #(int)::set(null,"*","PORT_1141_COUNT",port_count[1141]);
       uvm_config_db #(int)::set(null,"*","PORT_1142_COUNT",port_count[1142]);
       uvm_config_db #(int)::set(null,"*","PORT_1143_COUNT",port_count[1143]);
       uvm_config_db #(int)::set(null,"*","PORT_1144_COUNT",port_count[1144]);
       uvm_config_db #(int)::set(null,"*","PORT_1145_COUNT",port_count[1145]);
       uvm_config_db #(int)::set(null,"*","PORT_1146_COUNT",port_count[1146]);
       uvm_config_db #(int)::set(null,"*","PORT_1147_COUNT",port_count[1147]);
       uvm_config_db #(int)::set(null,"*","PORT_1148_COUNT",port_count[1148]);
       uvm_config_db #(int)::set(null,"*","PORT_1149_COUNT",port_count[1149]);
       uvm_config_db #(int)::set(null,"*","PORT_1150_COUNT",port_count[1150]);
       uvm_config_db #(int)::set(null,"*","PORT_1151_COUNT",port_count[1151]);
       uvm_config_db #(int)::set(null,"*","PORT_1152_COUNT",port_count[1152]);
       uvm_config_db #(int)::set(null,"*","PORT_1153_COUNT",port_count[1153]);
       uvm_config_db #(int)::set(null,"*","PORT_1154_COUNT",port_count[1154]);
       uvm_config_db #(int)::set(null,"*","PORT_1155_COUNT",port_count[1155]);
       uvm_config_db #(int)::set(null,"*","PORT_1156_COUNT",port_count[1156]);
       uvm_config_db #(int)::set(null,"*","PORT_1157_COUNT",port_count[1157]);
       uvm_config_db #(int)::set(null,"*","PORT_1158_COUNT",port_count[1158]);
       uvm_config_db #(int)::set(null,"*","PORT_1159_COUNT",port_count[1159]);
       uvm_config_db #(int)::set(null,"*","PORT_1160_COUNT",port_count[1160]);
       uvm_config_db #(int)::set(null,"*","PORT_1161_COUNT",port_count[1161]);
       uvm_config_db #(int)::set(null,"*","PORT_1162_COUNT",port_count[1162]);
       uvm_config_db #(int)::set(null,"*","PORT_1163_COUNT",port_count[1163]);
       uvm_config_db #(int)::set(null,"*","PORT_1164_COUNT",port_count[1164]);
       uvm_config_db #(int)::set(null,"*","PORT_1165_COUNT",port_count[1165]);
       uvm_config_db #(int)::set(null,"*","PORT_1166_COUNT",port_count[1166]);
       uvm_config_db #(int)::set(null,"*","PORT_1167_COUNT",port_count[1167]);
       uvm_config_db #(int)::set(null,"*","PORT_1168_COUNT",port_count[1168]);
       uvm_config_db #(int)::set(null,"*","PORT_1169_COUNT",port_count[1169]);
       uvm_config_db #(int)::set(null,"*","PORT_1170_COUNT",port_count[1170]);
       uvm_config_db #(int)::set(null,"*","PORT_1171_COUNT",port_count[1171]);
       uvm_config_db #(int)::set(null,"*","PORT_1172_COUNT",port_count[1172]);
       uvm_config_db #(int)::set(null,"*","PORT_1173_COUNT",port_count[1173]);
       uvm_config_db #(int)::set(null,"*","PORT_1174_COUNT",port_count[1174]);
       uvm_config_db #(int)::set(null,"*","PORT_1175_COUNT",port_count[1175]);
       uvm_config_db #(int)::set(null,"*","PORT_1176_COUNT",port_count[1176]);
       uvm_config_db #(int)::set(null,"*","PORT_1177_COUNT",port_count[1177]);
       uvm_config_db #(int)::set(null,"*","PORT_1178_COUNT",port_count[1178]);
       uvm_config_db #(int)::set(null,"*","PORT_1179_COUNT",port_count[1179]);
       uvm_config_db #(int)::set(null,"*","PORT_1180_COUNT",port_count[1180]);
       uvm_config_db #(int)::set(null,"*","PORT_1181_COUNT",port_count[1181]);
       uvm_config_db #(int)::set(null,"*","PORT_1182_COUNT",port_count[1182]);
       uvm_config_db #(int)::set(null,"*","PORT_1183_COUNT",port_count[1183]);
       uvm_config_db #(int)::set(null,"*","PORT_1184_COUNT",port_count[1184]);
       uvm_config_db #(int)::set(null,"*","PORT_1185_COUNT",port_count[1185]);
       uvm_config_db #(int)::set(null,"*","PORT_1186_COUNT",port_count[1186]);
       uvm_config_db #(int)::set(null,"*","PORT_1187_COUNT",port_count[1187]);
       uvm_config_db #(int)::set(null,"*","PORT_1188_COUNT",port_count[1188]);
       uvm_config_db #(int)::set(null,"*","PORT_1189_COUNT",port_count[1189]);
       uvm_config_db #(int)::set(null,"*","PORT_1190_COUNT",port_count[1190]);
       uvm_config_db #(int)::set(null,"*","PORT_1191_COUNT",port_count[1191]);
       uvm_config_db #(int)::set(null,"*","PORT_1192_COUNT",port_count[1192]);
       uvm_config_db #(int)::set(null,"*","PORT_1193_COUNT",port_count[1193]);
       uvm_config_db #(int)::set(null,"*","PORT_1194_COUNT",port_count[1194]);
       uvm_config_db #(int)::set(null,"*","PORT_1195_COUNT",port_count[1195]);
       uvm_config_db #(int)::set(null,"*","PORT_1196_COUNT",port_count[1196]);
       uvm_config_db #(int)::set(null,"*","PORT_1197_COUNT",port_count[1197]);
       uvm_config_db #(int)::set(null,"*","PORT_1198_COUNT",port_count[1198]);
       uvm_config_db #(int)::set(null,"*","PORT_1199_COUNT",port_count[1199]);
       uvm_config_db #(int)::set(null,"*","PORT_1200_COUNT",port_count[1200]);
       uvm_config_db #(int)::set(null,"*","PORT_1201_COUNT",port_count[1201]);
       uvm_config_db #(int)::set(null,"*","PORT_1202_COUNT",port_count[1202]);
       uvm_config_db #(int)::set(null,"*","PORT_1203_COUNT",port_count[1203]);
       uvm_config_db #(int)::set(null,"*","PORT_1204_COUNT",port_count[1204]);
       uvm_config_db #(int)::set(null,"*","PORT_1205_COUNT",port_count[1205]);
       uvm_config_db #(int)::set(null,"*","PORT_1206_COUNT",port_count[1206]);
       uvm_config_db #(int)::set(null,"*","PORT_1207_COUNT",port_count[1207]);
       uvm_config_db #(int)::set(null,"*","PORT_1208_COUNT",port_count[1208]);
       uvm_config_db #(int)::set(null,"*","PORT_1209_COUNT",port_count[1209]);
       uvm_config_db #(int)::set(null,"*","PORT_1210_COUNT",port_count[1210]);
       uvm_config_db #(int)::set(null,"*","PORT_1211_COUNT",port_count[1211]);
       uvm_config_db #(int)::set(null,"*","PORT_1212_COUNT",port_count[1212]);
       uvm_config_db #(int)::set(null,"*","PORT_1213_COUNT",port_count[1213]);
       uvm_config_db #(int)::set(null,"*","PORT_1214_COUNT",port_count[1214]);
       uvm_config_db #(int)::set(null,"*","PORT_1215_COUNT",port_count[1215]);
       uvm_config_db #(int)::set(null,"*","PORT_1216_COUNT",port_count[1216]);
       uvm_config_db #(int)::set(null,"*","PORT_1217_COUNT",port_count[1217]);
       uvm_config_db #(int)::set(null,"*","PORT_1218_COUNT",port_count[1218]);
       uvm_config_db #(int)::set(null,"*","PORT_1219_COUNT",port_count[1219]);
       uvm_config_db #(int)::set(null,"*","PORT_1220_COUNT",port_count[1220]);
       uvm_config_db #(int)::set(null,"*","PORT_1221_COUNT",port_count[1221]);
       uvm_config_db #(int)::set(null,"*","PORT_1222_COUNT",port_count[1222]);
       uvm_config_db #(int)::set(null,"*","PORT_1223_COUNT",port_count[1223]);
       uvm_config_db #(int)::set(null,"*","PORT_1224_COUNT",port_count[1224]);
       uvm_config_db #(int)::set(null,"*","PORT_1225_COUNT",port_count[1225]);
       uvm_config_db #(int)::set(null,"*","PORT_1226_COUNT",port_count[1226]);
       uvm_config_db #(int)::set(null,"*","PORT_1227_COUNT",port_count[1227]);
       uvm_config_db #(int)::set(null,"*","PORT_1228_COUNT",port_count[1228]);
       uvm_config_db #(int)::set(null,"*","PORT_1229_COUNT",port_count[1229]);
       uvm_config_db #(int)::set(null,"*","PORT_1230_COUNT",port_count[1230]);
       uvm_config_db #(int)::set(null,"*","PORT_1231_COUNT",port_count[1231]);
       uvm_config_db #(int)::set(null,"*","PORT_1232_COUNT",port_count[1232]);
       uvm_config_db #(int)::set(null,"*","PORT_1233_COUNT",port_count[1233]);
       uvm_config_db #(int)::set(null,"*","PORT_1234_COUNT",port_count[1234]);
       uvm_config_db #(int)::set(null,"*","PORT_1235_COUNT",port_count[1235]);
       uvm_config_db #(int)::set(null,"*","PORT_1236_COUNT",port_count[1236]);
       uvm_config_db #(int)::set(null,"*","PORT_1237_COUNT",port_count[1237]);
       uvm_config_db #(int)::set(null,"*","PORT_1238_COUNT",port_count[1238]);
       uvm_config_db #(int)::set(null,"*","PORT_1239_COUNT",port_count[1239]);
       uvm_config_db #(int)::set(null,"*","PORT_1240_COUNT",port_count[1240]);
       uvm_config_db #(int)::set(null,"*","PORT_1241_COUNT",port_count[1241]);
       uvm_config_db #(int)::set(null,"*","PORT_1242_COUNT",port_count[1242]);
       uvm_config_db #(int)::set(null,"*","PORT_1243_COUNT",port_count[1243]);
       uvm_config_db #(int)::set(null,"*","PORT_1244_COUNT",port_count[1244]);
       uvm_config_db #(int)::set(null,"*","PORT_1245_COUNT",port_count[1245]);
       uvm_config_db #(int)::set(null,"*","PORT_1246_COUNT",port_count[1246]);
       uvm_config_db #(int)::set(null,"*","PORT_1247_COUNT",port_count[1247]);
       uvm_config_db #(int)::set(null,"*","PORT_1248_COUNT",port_count[1248]);
       uvm_config_db #(int)::set(null,"*","PORT_1249_COUNT",port_count[1249]);
       uvm_config_db #(int)::set(null,"*","PORT_1250_COUNT",port_count[1250]);
       uvm_config_db #(int)::set(null,"*","PORT_1251_COUNT",port_count[1251]);
       uvm_config_db #(int)::set(null,"*","PORT_1252_COUNT",port_count[1252]);
       uvm_config_db #(int)::set(null,"*","PORT_1253_COUNT",port_count[1253]);
       uvm_config_db #(int)::set(null,"*","PORT_1254_COUNT",port_count[1254]);
       uvm_config_db #(int)::set(null,"*","PORT_1255_COUNT",port_count[1255]);
       uvm_config_db #(int)::set(null,"*","PORT_1256_COUNT",port_count[1256]);
       uvm_config_db #(int)::set(null,"*","PORT_1257_COUNT",port_count[1257]);
       uvm_config_db #(int)::set(null,"*","PORT_1258_COUNT",port_count[1258]);
       uvm_config_db #(int)::set(null,"*","PORT_1259_COUNT",port_count[1259]);
       uvm_config_db #(int)::set(null,"*","PORT_1260_COUNT",port_count[1260]);
       uvm_config_db #(int)::set(null,"*","PORT_1261_COUNT",port_count[1261]);
       uvm_config_db #(int)::set(null,"*","PORT_1262_COUNT",port_count[1262]);
       uvm_config_db #(int)::set(null,"*","PORT_1263_COUNT",port_count[1263]);
       uvm_config_db #(int)::set(null,"*","PORT_1264_COUNT",port_count[1264]);
       uvm_config_db #(int)::set(null,"*","PORT_1265_COUNT",port_count[1265]);
       uvm_config_db #(int)::set(null,"*","PORT_1266_COUNT",port_count[1266]);
       uvm_config_db #(int)::set(null,"*","PORT_1267_COUNT",port_count[1267]);
       uvm_config_db #(int)::set(null,"*","PORT_1268_COUNT",port_count[1268]);
       uvm_config_db #(int)::set(null,"*","PORT_1269_COUNT",port_count[1269]);
       uvm_config_db #(int)::set(null,"*","PORT_1270_COUNT",port_count[1270]);
       uvm_config_db #(int)::set(null,"*","PORT_1271_COUNT",port_count[1271]);
       uvm_config_db #(int)::set(null,"*","PORT_1272_COUNT",port_count[1272]);
       uvm_config_db #(int)::set(null,"*","PORT_1273_COUNT",port_count[1273]);
       uvm_config_db #(int)::set(null,"*","PORT_1274_COUNT",port_count[1274]);
       uvm_config_db #(int)::set(null,"*","PORT_1275_COUNT",port_count[1275]);
       uvm_config_db #(int)::set(null,"*","PORT_1276_COUNT",port_count[1276]);
       uvm_config_db #(int)::set(null,"*","PORT_1277_COUNT",port_count[1277]);
       uvm_config_db #(int)::set(null,"*","PORT_1278_COUNT",port_count[1278]);
       uvm_config_db #(int)::set(null,"*","PORT_1279_COUNT",port_count[1279]);
       uvm_config_db #(int)::set(null,"*","PORT_1280_COUNT",port_count[1280]);
       uvm_config_db #(int)::set(null,"*","PORT_1281_COUNT",port_count[1281]);
       uvm_config_db #(int)::set(null,"*","PORT_1282_COUNT",port_count[1282]);
       uvm_config_db #(int)::set(null,"*","PORT_1283_COUNT",port_count[1283]);
       uvm_config_db #(int)::set(null,"*","PORT_1284_COUNT",port_count[1284]);
       uvm_config_db #(int)::set(null,"*","PORT_1285_COUNT",port_count[1285]);
       uvm_config_db #(int)::set(null,"*","PORT_1286_COUNT",port_count[1286]);
       uvm_config_db #(int)::set(null,"*","PORT_1287_COUNT",port_count[1287]);
       uvm_config_db #(int)::set(null,"*","PORT_1288_COUNT",port_count[1288]);
       uvm_config_db #(int)::set(null,"*","PORT_1289_COUNT",port_count[1289]);
       uvm_config_db #(int)::set(null,"*","PORT_1290_COUNT",port_count[1290]);
       uvm_config_db #(int)::set(null,"*","PORT_1291_COUNT",port_count[1291]);
       uvm_config_db #(int)::set(null,"*","PORT_1292_COUNT",port_count[1292]);
       uvm_config_db #(int)::set(null,"*","PORT_1293_COUNT",port_count[1293]);
       uvm_config_db #(int)::set(null,"*","PORT_1294_COUNT",port_count[1294]);
       uvm_config_db #(int)::set(null,"*","PORT_1295_COUNT",port_count[1295]);
       uvm_config_db #(int)::set(null,"*","PORT_1296_COUNT",port_count[1296]);
       uvm_config_db #(int)::set(null,"*","PORT_1297_COUNT",port_count[1297]);
       uvm_config_db #(int)::set(null,"*","PORT_1298_COUNT",port_count[1298]);
       uvm_config_db #(int)::set(null,"*","PORT_1299_COUNT",port_count[1299]);
       uvm_config_db #(int)::set(null,"*","PORT_1300_COUNT",port_count[1300]);
       uvm_config_db #(int)::set(null,"*","PORT_1301_COUNT",port_count[1301]);
       uvm_config_db #(int)::set(null,"*","PORT_1302_COUNT",port_count[1302]);
       uvm_config_db #(int)::set(null,"*","PORT_1303_COUNT",port_count[1303]);
       uvm_config_db #(int)::set(null,"*","PORT_1304_COUNT",port_count[1304]);
       uvm_config_db #(int)::set(null,"*","PORT_1305_COUNT",port_count[1305]);
       uvm_config_db #(int)::set(null,"*","PORT_1306_COUNT",port_count[1306]);
       uvm_config_db #(int)::set(null,"*","PORT_1307_COUNT",port_count[1307]);
       uvm_config_db #(int)::set(null,"*","PORT_1308_COUNT",port_count[1308]);
       uvm_config_db #(int)::set(null,"*","PORT_1309_COUNT",port_count[1309]);
       uvm_config_db #(int)::set(null,"*","PORT_1310_COUNT",port_count[1310]);
       uvm_config_db #(int)::set(null,"*","PORT_1311_COUNT",port_count[1311]);
       uvm_config_db #(int)::set(null,"*","PORT_1312_COUNT",port_count[1312]);
       uvm_config_db #(int)::set(null,"*","PORT_1313_COUNT",port_count[1313]);
       uvm_config_db #(int)::set(null,"*","PORT_1314_COUNT",port_count[1314]);
       uvm_config_db #(int)::set(null,"*","PORT_1315_COUNT",port_count[1315]);
       uvm_config_db #(int)::set(null,"*","PORT_1316_COUNT",port_count[1316]);
       uvm_config_db #(int)::set(null,"*","PORT_1317_COUNT",port_count[1317]);
       uvm_config_db #(int)::set(null,"*","PORT_1318_COUNT",port_count[1318]);
       uvm_config_db #(int)::set(null,"*","PORT_1319_COUNT",port_count[1319]);
       uvm_config_db #(int)::set(null,"*","PORT_1320_COUNT",port_count[1320]);
       uvm_config_db #(int)::set(null,"*","PORT_1321_COUNT",port_count[1321]);
       uvm_config_db #(int)::set(null,"*","PORT_1322_COUNT",port_count[1322]);
       uvm_config_db #(int)::set(null,"*","PORT_1323_COUNT",port_count[1323]);
       uvm_config_db #(int)::set(null,"*","PORT_1324_COUNT",port_count[1324]);
       uvm_config_db #(int)::set(null,"*","PORT_1325_COUNT",port_count[1325]);
       uvm_config_db #(int)::set(null,"*","PORT_1326_COUNT",port_count[1326]);
       uvm_config_db #(int)::set(null,"*","PORT_1327_COUNT",port_count[1327]);
       uvm_config_db #(int)::set(null,"*","PORT_1328_COUNT",port_count[1328]);
       uvm_config_db #(int)::set(null,"*","PORT_1329_COUNT",port_count[1329]);
       uvm_config_db #(int)::set(null,"*","PORT_1330_COUNT",port_count[1330]);
       uvm_config_db #(int)::set(null,"*","PORT_1331_COUNT",port_count[1331]);
       uvm_config_db #(int)::set(null,"*","PORT_1332_COUNT",port_count[1332]);
       uvm_config_db #(int)::set(null,"*","PORT_1333_COUNT",port_count[1333]);
       uvm_config_db #(int)::set(null,"*","PORT_1334_COUNT",port_count[1334]);
       uvm_config_db #(int)::set(null,"*","PORT_1335_COUNT",port_count[1335]);
       uvm_config_db #(int)::set(null,"*","PORT_1336_COUNT",port_count[1336]);
       uvm_config_db #(int)::set(null,"*","PORT_1337_COUNT",port_count[1337]);
       uvm_config_db #(int)::set(null,"*","PORT_1338_COUNT",port_count[1338]);
       uvm_config_db #(int)::set(null,"*","PORT_1339_COUNT",port_count[1339]);
       uvm_config_db #(int)::set(null,"*","PORT_1340_COUNT",port_count[1340]);
       uvm_config_db #(int)::set(null,"*","PORT_1341_COUNT",port_count[1341]);
       uvm_config_db #(int)::set(null,"*","PORT_1342_COUNT",port_count[1342]);
       uvm_config_db #(int)::set(null,"*","PORT_1343_COUNT",port_count[1343]);
       uvm_config_db #(int)::set(null,"*","PORT_1344_COUNT",port_count[1344]);
       uvm_config_db #(int)::set(null,"*","PORT_1345_COUNT",port_count[1345]);
       uvm_config_db #(int)::set(null,"*","PORT_1346_COUNT",port_count[1346]);
       uvm_config_db #(int)::set(null,"*","PORT_1347_COUNT",port_count[1347]);
       uvm_config_db #(int)::set(null,"*","PORT_1348_COUNT",port_count[1348]);
       uvm_config_db #(int)::set(null,"*","PORT_1349_COUNT",port_count[1349]);
       uvm_config_db #(int)::set(null,"*","PORT_1350_COUNT",port_count[1350]);
       uvm_config_db #(int)::set(null,"*","PORT_1351_COUNT",port_count[1351]);
       uvm_config_db #(int)::set(null,"*","PORT_1352_COUNT",port_count[1352]);
       uvm_config_db #(int)::set(null,"*","PORT_1353_COUNT",port_count[1353]);
       uvm_config_db #(int)::set(null,"*","PORT_1354_COUNT",port_count[1354]);
       uvm_config_db #(int)::set(null,"*","PORT_1355_COUNT",port_count[1355]);
       uvm_config_db #(int)::set(null,"*","PORT_1356_COUNT",port_count[1356]);
       uvm_config_db #(int)::set(null,"*","PORT_1357_COUNT",port_count[1357]);
       uvm_config_db #(int)::set(null,"*","PORT_1358_COUNT",port_count[1358]);
       uvm_config_db #(int)::set(null,"*","PORT_1359_COUNT",port_count[1359]);
       uvm_config_db #(int)::set(null,"*","PORT_1360_COUNT",port_count[1360]);
       uvm_config_db #(int)::set(null,"*","PORT_1361_COUNT",port_count[1361]);
       uvm_config_db #(int)::set(null,"*","PORT_1362_COUNT",port_count[1362]);
       uvm_config_db #(int)::set(null,"*","PORT_1363_COUNT",port_count[1363]);
       uvm_config_db #(int)::set(null,"*","PORT_1364_COUNT",port_count[1364]);
       uvm_config_db #(int)::set(null,"*","PORT_1365_COUNT",port_count[1365]);
       uvm_config_db #(int)::set(null,"*","PORT_1366_COUNT",port_count[1366]);
       uvm_config_db #(int)::set(null,"*","PORT_1367_COUNT",port_count[1367]);
       uvm_config_db #(int)::set(null,"*","PORT_1368_COUNT",port_count[1368]);
       uvm_config_db #(int)::set(null,"*","PORT_1369_COUNT",port_count[1369]);
       uvm_config_db #(int)::set(null,"*","PORT_1370_COUNT",port_count[1370]);
       uvm_config_db #(int)::set(null,"*","PORT_1371_COUNT",port_count[1371]);
       uvm_config_db #(int)::set(null,"*","PORT_1372_COUNT",port_count[1372]);
       uvm_config_db #(int)::set(null,"*","PORT_1373_COUNT",port_count[1373]);
       uvm_config_db #(int)::set(null,"*","PORT_1374_COUNT",port_count[1374]);
       uvm_config_db #(int)::set(null,"*","PORT_1375_COUNT",port_count[1375]);
       uvm_config_db #(int)::set(null,"*","PORT_1376_COUNT",port_count[1376]);
       uvm_config_db #(int)::set(null,"*","PORT_1377_COUNT",port_count[1377]);
       uvm_config_db #(int)::set(null,"*","PORT_1378_COUNT",port_count[1378]);
       uvm_config_db #(int)::set(null,"*","PORT_1379_COUNT",port_count[1379]);
       uvm_config_db #(int)::set(null,"*","PORT_1380_COUNT",port_count[1380]);
       uvm_config_db #(int)::set(null,"*","PORT_1381_COUNT",port_count[1381]);
       uvm_config_db #(int)::set(null,"*","PORT_1382_COUNT",port_count[1382]);
       uvm_config_db #(int)::set(null,"*","PORT_1383_COUNT",port_count[1383]);
       uvm_config_db #(int)::set(null,"*","PORT_1384_COUNT",port_count[1384]);
       uvm_config_db #(int)::set(null,"*","PORT_1385_COUNT",port_count[1385]);
       uvm_config_db #(int)::set(null,"*","PORT_1386_COUNT",port_count[1386]);
       uvm_config_db #(int)::set(null,"*","PORT_1387_COUNT",port_count[1387]);
       uvm_config_db #(int)::set(null,"*","PORT_1388_COUNT",port_count[1388]);
       uvm_config_db #(int)::set(null,"*","PORT_1389_COUNT",port_count[1389]);
       uvm_config_db #(int)::set(null,"*","PORT_1390_COUNT",port_count[1390]);
       uvm_config_db #(int)::set(null,"*","PORT_1391_COUNT",port_count[1391]);
       uvm_config_db #(int)::set(null,"*","PORT_1392_COUNT",port_count[1392]);
       uvm_config_db #(int)::set(null,"*","PORT_1393_COUNT",port_count[1393]);
       uvm_config_db #(int)::set(null,"*","PORT_1394_COUNT",port_count[1394]);
       uvm_config_db #(int)::set(null,"*","PORT_1395_COUNT",port_count[1395]);
       uvm_config_db #(int)::set(null,"*","PORT_1396_COUNT",port_count[1396]);
       uvm_config_db #(int)::set(null,"*","PORT_1397_COUNT",port_count[1397]);
       uvm_config_db #(int)::set(null,"*","PORT_1398_COUNT",port_count[1398]);
       uvm_config_db #(int)::set(null,"*","PORT_1399_COUNT",port_count[1399]);
       uvm_config_db #(int)::set(null,"*","PORT_1400_COUNT",port_count[1400]);
       uvm_config_db #(int)::set(null,"*","PORT_1401_COUNT",port_count[1401]);
       uvm_config_db #(int)::set(null,"*","PORT_1402_COUNT",port_count[1402]);
       uvm_config_db #(int)::set(null,"*","PORT_1403_COUNT",port_count[1403]);
       uvm_config_db #(int)::set(null,"*","PORT_1404_COUNT",port_count[1404]);
       uvm_config_db #(int)::set(null,"*","PORT_1405_COUNT",port_count[1405]);
       uvm_config_db #(int)::set(null,"*","PORT_1406_COUNT",port_count[1406]);
       uvm_config_db #(int)::set(null,"*","PORT_1407_COUNT",port_count[1407]);
       uvm_config_db #(int)::set(null,"*","PORT_1408_COUNT",port_count[1408]);
       uvm_config_db #(int)::set(null,"*","PORT_1409_COUNT",port_count[1409]);
       uvm_config_db #(int)::set(null,"*","PORT_1410_COUNT",port_count[1410]);
       uvm_config_db #(int)::set(null,"*","PORT_1411_COUNT",port_count[1411]);
       uvm_config_db #(int)::set(null,"*","PORT_1412_COUNT",port_count[1412]);
       uvm_config_db #(int)::set(null,"*","PORT_1413_COUNT",port_count[1413]);
       uvm_config_db #(int)::set(null,"*","PORT_1414_COUNT",port_count[1414]);
       uvm_config_db #(int)::set(null,"*","PORT_1415_COUNT",port_count[1415]);
       uvm_config_db #(int)::set(null,"*","PORT_1416_COUNT",port_count[1416]);
       uvm_config_db #(int)::set(null,"*","PORT_1417_COUNT",port_count[1417]);
       uvm_config_db #(int)::set(null,"*","PORT_1418_COUNT",port_count[1418]);
       uvm_config_db #(int)::set(null,"*","PORT_1419_COUNT",port_count[1419]);
       uvm_config_db #(int)::set(null,"*","PORT_1420_COUNT",port_count[1420]);
       uvm_config_db #(int)::set(null,"*","PORT_1421_COUNT",port_count[1421]);
       uvm_config_db #(int)::set(null,"*","PORT_1422_COUNT",port_count[1422]);
       uvm_config_db #(int)::set(null,"*","PORT_1423_COUNT",port_count[1423]);
       uvm_config_db #(int)::set(null,"*","PORT_1424_COUNT",port_count[1424]);
       uvm_config_db #(int)::set(null,"*","PORT_1425_COUNT",port_count[1425]);
       uvm_config_db #(int)::set(null,"*","PORT_1426_COUNT",port_count[1426]);
       uvm_config_db #(int)::set(null,"*","PORT_1427_COUNT",port_count[1427]);
       uvm_config_db #(int)::set(null,"*","PORT_1428_COUNT",port_count[1428]);
       uvm_config_db #(int)::set(null,"*","PORT_1429_COUNT",port_count[1429]);
       uvm_config_db #(int)::set(null,"*","PORT_1430_COUNT",port_count[1430]);
       uvm_config_db #(int)::set(null,"*","PORT_1431_COUNT",port_count[1431]);
       uvm_config_db #(int)::set(null,"*","PORT_1432_COUNT",port_count[1432]);
       uvm_config_db #(int)::set(null,"*","PORT_1433_COUNT",port_count[1433]);
       uvm_config_db #(int)::set(null,"*","PORT_1434_COUNT",port_count[1434]);
       uvm_config_db #(int)::set(null,"*","PORT_1435_COUNT",port_count[1435]);
       uvm_config_db #(int)::set(null,"*","PORT_1436_COUNT",port_count[1436]);
       uvm_config_db #(int)::set(null,"*","PORT_1437_COUNT",port_count[1437]);
       uvm_config_db #(int)::set(null,"*","PORT_1438_COUNT",port_count[1438]);
       uvm_config_db #(int)::set(null,"*","PORT_1439_COUNT",port_count[1439]);
       uvm_config_db #(int)::set(null,"*","PORT_1440_COUNT",port_count[1440]);
       uvm_config_db #(int)::set(null,"*","PORT_1441_COUNT",port_count[1441]);
       uvm_config_db #(int)::set(null,"*","PORT_1442_COUNT",port_count[1442]);
       uvm_config_db #(int)::set(null,"*","PORT_1443_COUNT",port_count[1443]);
       uvm_config_db #(int)::set(null,"*","PORT_1444_COUNT",port_count[1444]);
       uvm_config_db #(int)::set(null,"*","PORT_1445_COUNT",port_count[1445]);
       uvm_config_db #(int)::set(null,"*","PORT_1446_COUNT",port_count[1446]);
       uvm_config_db #(int)::set(null,"*","PORT_1447_COUNT",port_count[1447]);
       uvm_config_db #(int)::set(null,"*","PORT_1448_COUNT",port_count[1448]);
       uvm_config_db #(int)::set(null,"*","PORT_1449_COUNT",port_count[1449]);
       uvm_config_db #(int)::set(null,"*","PORT_1450_COUNT",port_count[1450]);
       uvm_config_db #(int)::set(null,"*","PORT_1451_COUNT",port_count[1451]);
       uvm_config_db #(int)::set(null,"*","PORT_1452_COUNT",port_count[1452]);
       uvm_config_db #(int)::set(null,"*","PORT_1453_COUNT",port_count[1453]);
       uvm_config_db #(int)::set(null,"*","PORT_1454_COUNT",port_count[1454]);
       uvm_config_db #(int)::set(null,"*","PORT_1455_COUNT",port_count[1455]);
       uvm_config_db #(int)::set(null,"*","PORT_1456_COUNT",port_count[1456]);
       uvm_config_db #(int)::set(null,"*","PORT_1457_COUNT",port_count[1457]);
       uvm_config_db #(int)::set(null,"*","PORT_1458_COUNT",port_count[1458]);
       uvm_config_db #(int)::set(null,"*","PORT_1459_COUNT",port_count[1459]);
       uvm_config_db #(int)::set(null,"*","PORT_1460_COUNT",port_count[1460]);
       uvm_config_db #(int)::set(null,"*","PORT_1461_COUNT",port_count[1461]);
       uvm_config_db #(int)::set(null,"*","PORT_1462_COUNT",port_count[1462]);
       uvm_config_db #(int)::set(null,"*","PORT_1463_COUNT",port_count[1463]);
       uvm_config_db #(int)::set(null,"*","PORT_1464_COUNT",port_count[1464]);
       uvm_config_db #(int)::set(null,"*","PORT_1465_COUNT",port_count[1465]);
       uvm_config_db #(int)::set(null,"*","PORT_1466_COUNT",port_count[1466]);
       uvm_config_db #(int)::set(null,"*","PORT_1467_COUNT",port_count[1467]);
       uvm_config_db #(int)::set(null,"*","PORT_1468_COUNT",port_count[1468]);
       uvm_config_db #(int)::set(null,"*","PORT_1469_COUNT",port_count[1469]);
       uvm_config_db #(int)::set(null,"*","PORT_1470_COUNT",port_count[1470]);
       uvm_config_db #(int)::set(null,"*","PORT_1471_COUNT",port_count[1471]);
       uvm_config_db #(int)::set(null,"*","PORT_1472_COUNT",port_count[1472]);
       uvm_config_db #(int)::set(null,"*","PORT_1473_COUNT",port_count[1473]);
       uvm_config_db #(int)::set(null,"*","PORT_1474_COUNT",port_count[1474]);
       uvm_config_db #(int)::set(null,"*","PORT_1475_COUNT",port_count[1475]);
       uvm_config_db #(int)::set(null,"*","PORT_1476_COUNT",port_count[1476]);
       uvm_config_db #(int)::set(null,"*","PORT_1477_COUNT",port_count[1477]);
       uvm_config_db #(int)::set(null,"*","PORT_1478_COUNT",port_count[1478]);
       uvm_config_db #(int)::set(null,"*","PORT_1479_COUNT",port_count[1479]);
       uvm_config_db #(int)::set(null,"*","PORT_1480_COUNT",port_count[1480]);
       uvm_config_db #(int)::set(null,"*","PORT_1481_COUNT",port_count[1481]);
       uvm_config_db #(int)::set(null,"*","PORT_1482_COUNT",port_count[1482]);
       uvm_config_db #(int)::set(null,"*","PORT_1483_COUNT",port_count[1483]);
       uvm_config_db #(int)::set(null,"*","PORT_1484_COUNT",port_count[1484]);
       uvm_config_db #(int)::set(null,"*","PORT_1485_COUNT",port_count[1485]);
       uvm_config_db #(int)::set(null,"*","PORT_1486_COUNT",port_count[1486]);
       uvm_config_db #(int)::set(null,"*","PORT_1487_COUNT",port_count[1487]);
       uvm_config_db #(int)::set(null,"*","PORT_1488_COUNT",port_count[1488]);
       uvm_config_db #(int)::set(null,"*","PORT_1489_COUNT",port_count[1489]);
       uvm_config_db #(int)::set(null,"*","PORT_1490_COUNT",port_count[1490]);
       uvm_config_db #(int)::set(null,"*","PORT_1491_COUNT",port_count[1491]);
       uvm_config_db #(int)::set(null,"*","PORT_1492_COUNT",port_count[1492]);
       uvm_config_db #(int)::set(null,"*","PORT_1493_COUNT",port_count[1493]);
       uvm_config_db #(int)::set(null,"*","PORT_1494_COUNT",port_count[1494]);
       uvm_config_db #(int)::set(null,"*","PORT_1495_COUNT",port_count[1495]);
       uvm_config_db #(int)::set(null,"*","PORT_1496_COUNT",port_count[1496]);
       uvm_config_db #(int)::set(null,"*","PORT_1497_COUNT",port_count[1497]);
       uvm_config_db #(int)::set(null,"*","PORT_1498_COUNT",port_count[1498]);
       uvm_config_db #(int)::set(null,"*","PORT_1499_COUNT",port_count[1499]);
       uvm_config_db #(int)::set(null,"*","PORT_1500_COUNT",port_count[1500]);
       uvm_config_db #(int)::set(null,"*","PORT_1501_COUNT",port_count[1501]);
       uvm_config_db #(int)::set(null,"*","PORT_1502_COUNT",port_count[1502]);
       uvm_config_db #(int)::set(null,"*","PORT_1503_COUNT",port_count[1503]);
       uvm_config_db #(int)::set(null,"*","PORT_1504_COUNT",port_count[1504]);
       uvm_config_db #(int)::set(null,"*","PORT_1505_COUNT",port_count[1505]);
       uvm_config_db #(int)::set(null,"*","PORT_1506_COUNT",port_count[1506]);
       uvm_config_db #(int)::set(null,"*","PORT_1507_COUNT",port_count[1507]);
       uvm_config_db #(int)::set(null,"*","PORT_1508_COUNT",port_count[1508]);
       uvm_config_db #(int)::set(null,"*","PORT_1509_COUNT",port_count[1509]);
       uvm_config_db #(int)::set(null,"*","PORT_1510_COUNT",port_count[1510]);
       uvm_config_db #(int)::set(null,"*","PORT_1511_COUNT",port_count[1511]);
       uvm_config_db #(int)::set(null,"*","PORT_1512_COUNT",port_count[1512]);
       uvm_config_db #(int)::set(null,"*","PORT_1513_COUNT",port_count[1513]);
       uvm_config_db #(int)::set(null,"*","PORT_1514_COUNT",port_count[1514]);
       uvm_config_db #(int)::set(null,"*","PORT_1515_COUNT",port_count[1515]);
       uvm_config_db #(int)::set(null,"*","PORT_1516_COUNT",port_count[1516]);
       uvm_config_db #(int)::set(null,"*","PORT_1517_COUNT",port_count[1517]);
       uvm_config_db #(int)::set(null,"*","PORT_1518_COUNT",port_count[1518]);
       uvm_config_db #(int)::set(null,"*","PORT_1519_COUNT",port_count[1519]);
       uvm_config_db #(int)::set(null,"*","PORT_1520_COUNT",port_count[1520]);
       uvm_config_db #(int)::set(null,"*","PORT_1521_COUNT",port_count[1521]);
       uvm_config_db #(int)::set(null,"*","PORT_1522_COUNT",port_count[1522]);
       uvm_config_db #(int)::set(null,"*","PORT_1523_COUNT",port_count[1523]);
       uvm_config_db #(int)::set(null,"*","PORT_1524_COUNT",port_count[1524]);
       uvm_config_db #(int)::set(null,"*","PORT_1525_COUNT",port_count[1525]);
       uvm_config_db #(int)::set(null,"*","PORT_1526_COUNT",port_count[1526]);
       uvm_config_db #(int)::set(null,"*","PORT_1527_COUNT",port_count[1527]);
       uvm_config_db #(int)::set(null,"*","PORT_1528_COUNT",port_count[1528]);
       uvm_config_db #(int)::set(null,"*","PORT_1529_COUNT",port_count[1529]);
       uvm_config_db #(int)::set(null,"*","PORT_1530_COUNT",port_count[1530]);
       uvm_config_db #(int)::set(null,"*","PORT_1531_COUNT",port_count[1531]);
       uvm_config_db #(int)::set(null,"*","PORT_1532_COUNT",port_count[1532]);
       uvm_config_db #(int)::set(null,"*","PORT_1533_COUNT",port_count[1533]);
       uvm_config_db #(int)::set(null,"*","PORT_1534_COUNT",port_count[1534]);
       uvm_config_db #(int)::set(null,"*","PORT_1535_COUNT",port_count[1535]);
       uvm_config_db #(int)::set(null,"*","PORT_1536_COUNT",port_count[1536]);
       uvm_config_db #(int)::set(null,"*","PORT_1537_COUNT",port_count[1537]);
       uvm_config_db #(int)::set(null,"*","PORT_1538_COUNT",port_count[1538]);
       uvm_config_db #(int)::set(null,"*","PORT_1539_COUNT",port_count[1539]);
       uvm_config_db #(int)::set(null,"*","PORT_1540_COUNT",port_count[1540]);
       uvm_config_db #(int)::set(null,"*","PORT_1541_COUNT",port_count[1541]);
       uvm_config_db #(int)::set(null,"*","PORT_1542_COUNT",port_count[1542]);
       uvm_config_db #(int)::set(null,"*","PORT_1543_COUNT",port_count[1543]);
       uvm_config_db #(int)::set(null,"*","PORT_1544_COUNT",port_count[1544]);
       uvm_config_db #(int)::set(null,"*","PORT_1545_COUNT",port_count[1545]);
       uvm_config_db #(int)::set(null,"*","PORT_1546_COUNT",port_count[1546]);
       uvm_config_db #(int)::set(null,"*","PORT_1547_COUNT",port_count[1547]);
       uvm_config_db #(int)::set(null,"*","PORT_1548_COUNT",port_count[1548]);
       uvm_config_db #(int)::set(null,"*","PORT_1549_COUNT",port_count[1549]);
       uvm_config_db #(int)::set(null,"*","PORT_1550_COUNT",port_count[1550]);
       uvm_config_db #(int)::set(null,"*","PORT_1551_COUNT",port_count[1551]);
       uvm_config_db #(int)::set(null,"*","PORT_1552_COUNT",port_count[1552]);
       uvm_config_db #(int)::set(null,"*","PORT_1553_COUNT",port_count[1553]);
       uvm_config_db #(int)::set(null,"*","PORT_1554_COUNT",port_count[1554]);
       uvm_config_db #(int)::set(null,"*","PORT_1555_COUNT",port_count[1555]);
       uvm_config_db #(int)::set(null,"*","PORT_1556_COUNT",port_count[1556]);
       uvm_config_db #(int)::set(null,"*","PORT_1557_COUNT",port_count[1557]);
       uvm_config_db #(int)::set(null,"*","PORT_1558_COUNT",port_count[1558]);
       uvm_config_db #(int)::set(null,"*","PORT_1559_COUNT",port_count[1559]);
       uvm_config_db #(int)::set(null,"*","PORT_1560_COUNT",port_count[1560]);
       uvm_config_db #(int)::set(null,"*","PORT_1561_COUNT",port_count[1561]);
       uvm_config_db #(int)::set(null,"*","PORT_1562_COUNT",port_count[1562]);
       uvm_config_db #(int)::set(null,"*","PORT_1563_COUNT",port_count[1563]);
       uvm_config_db #(int)::set(null,"*","PORT_1564_COUNT",port_count[1564]);
       uvm_config_db #(int)::set(null,"*","PORT_1565_COUNT",port_count[1565]);
       uvm_config_db #(int)::set(null,"*","PORT_1566_COUNT",port_count[1566]);
       uvm_config_db #(int)::set(null,"*","PORT_1567_COUNT",port_count[1567]);
       uvm_config_db #(int)::set(null,"*","PORT_1568_COUNT",port_count[1568]);
       uvm_config_db #(int)::set(null,"*","PORT_1569_COUNT",port_count[1569]);
       uvm_config_db #(int)::set(null,"*","PORT_1570_COUNT",port_count[1570]);
       uvm_config_db #(int)::set(null,"*","PORT_1571_COUNT",port_count[1571]);
       uvm_config_db #(int)::set(null,"*","PORT_1572_COUNT",port_count[1572]);
       uvm_config_db #(int)::set(null,"*","PORT_1573_COUNT",port_count[1573]);
       uvm_config_db #(int)::set(null,"*","PORT_1574_COUNT",port_count[1574]);
       uvm_config_db #(int)::set(null,"*","PORT_1575_COUNT",port_count[1575]);
       uvm_config_db #(int)::set(null,"*","PORT_1576_COUNT",port_count[1576]);
       uvm_config_db #(int)::set(null,"*","PORT_1577_COUNT",port_count[1577]);
       uvm_config_db #(int)::set(null,"*","PORT_1578_COUNT",port_count[1578]);
       uvm_config_db #(int)::set(null,"*","PORT_1579_COUNT",port_count[1579]);
       uvm_config_db #(int)::set(null,"*","PORT_1580_COUNT",port_count[1580]);
       uvm_config_db #(int)::set(null,"*","PORT_1581_COUNT",port_count[1581]);
       uvm_config_db #(int)::set(null,"*","PORT_1582_COUNT",port_count[1582]);
       uvm_config_db #(int)::set(null,"*","PORT_1583_COUNT",port_count[1583]);
       uvm_config_db #(int)::set(null,"*","PORT_1584_COUNT",port_count[1584]);
       uvm_config_db #(int)::set(null,"*","PORT_1585_COUNT",port_count[1585]);
       uvm_config_db #(int)::set(null,"*","PORT_1586_COUNT",port_count[1586]);
       uvm_config_db #(int)::set(null,"*","PORT_1587_COUNT",port_count[1587]);
       uvm_config_db #(int)::set(null,"*","PORT_1588_COUNT",port_count[1588]);
       uvm_config_db #(int)::set(null,"*","PORT_1589_COUNT",port_count[1589]);
       uvm_config_db #(int)::set(null,"*","PORT_1590_COUNT",port_count[1590]);
       uvm_config_db #(int)::set(null,"*","PORT_1591_COUNT",port_count[1591]);
       uvm_config_db #(int)::set(null,"*","PORT_1592_COUNT",port_count[1592]);
       uvm_config_db #(int)::set(null,"*","PORT_1593_COUNT",port_count[1593]);
       uvm_config_db #(int)::set(null,"*","PORT_1594_COUNT",port_count[1594]);
       uvm_config_db #(int)::set(null,"*","PORT_1595_COUNT",port_count[1595]);
       uvm_config_db #(int)::set(null,"*","PORT_1596_COUNT",port_count[1596]);
       uvm_config_db #(int)::set(null,"*","PORT_1597_COUNT",port_count[1597]);
       uvm_config_db #(int)::set(null,"*","PORT_1598_COUNT",port_count[1598]);
       uvm_config_db #(int)::set(null,"*","PORT_1599_COUNT",port_count[1599]);
       uvm_config_db #(int)::set(null,"*","PORT_1600_COUNT",port_count[1600]);
       uvm_config_db #(int)::set(null,"*","PORT_1601_COUNT",port_count[1601]);
       uvm_config_db #(int)::set(null,"*","PORT_1602_COUNT",port_count[1602]);
       uvm_config_db #(int)::set(null,"*","PORT_1603_COUNT",port_count[1603]);
       uvm_config_db #(int)::set(null,"*","PORT_1604_COUNT",port_count[1604]);
       uvm_config_db #(int)::set(null,"*","PORT_1605_COUNT",port_count[1605]);
       uvm_config_db #(int)::set(null,"*","PORT_1606_COUNT",port_count[1606]);
       uvm_config_db #(int)::set(null,"*","PORT_1607_COUNT",port_count[1607]);
       uvm_config_db #(int)::set(null,"*","PORT_1608_COUNT",port_count[1608]);
       uvm_config_db #(int)::set(null,"*","PORT_1609_COUNT",port_count[1609]);
       uvm_config_db #(int)::set(null,"*","PORT_1610_COUNT",port_count[1610]);
       uvm_config_db #(int)::set(null,"*","PORT_1611_COUNT",port_count[1611]);
       uvm_config_db #(int)::set(null,"*","PORT_1612_COUNT",port_count[1612]);
       uvm_config_db #(int)::set(null,"*","PORT_1613_COUNT",port_count[1613]);
       uvm_config_db #(int)::set(null,"*","PORT_1614_COUNT",port_count[1614]);
       uvm_config_db #(int)::set(null,"*","PORT_1615_COUNT",port_count[1615]);
       uvm_config_db #(int)::set(null,"*","PORT_1616_COUNT",port_count[1616]);
       uvm_config_db #(int)::set(null,"*","PORT_1617_COUNT",port_count[1617]);
       uvm_config_db #(int)::set(null,"*","PORT_1618_COUNT",port_count[1618]);
       uvm_config_db #(int)::set(null,"*","PORT_1619_COUNT",port_count[1619]);
       uvm_config_db #(int)::set(null,"*","PORT_1620_COUNT",port_count[1620]);
       uvm_config_db #(int)::set(null,"*","PORT_1621_COUNT",port_count[1621]);
       uvm_config_db #(int)::set(null,"*","PORT_1622_COUNT",port_count[1622]);
       uvm_config_db #(int)::set(null,"*","PORT_1623_COUNT",port_count[1623]);
       uvm_config_db #(int)::set(null,"*","PORT_1624_COUNT",port_count[1624]);
       uvm_config_db #(int)::set(null,"*","PORT_1625_COUNT",port_count[1625]);
       uvm_config_db #(int)::set(null,"*","PORT_1626_COUNT",port_count[1626]);
       uvm_config_db #(int)::set(null,"*","PORT_1627_COUNT",port_count[1627]);
       uvm_config_db #(int)::set(null,"*","PORT_1628_COUNT",port_count[1628]);
       uvm_config_db #(int)::set(null,"*","PORT_1629_COUNT",port_count[1629]);
       uvm_config_db #(int)::set(null,"*","PORT_1630_COUNT",port_count[1630]);
       uvm_config_db #(int)::set(null,"*","PORT_1631_COUNT",port_count[1631]);
       uvm_config_db #(int)::set(null,"*","PORT_1632_COUNT",port_count[1632]);
       uvm_config_db #(int)::set(null,"*","PORT_1633_COUNT",port_count[1633]);
       uvm_config_db #(int)::set(null,"*","PORT_1634_COUNT",port_count[1634]);
       uvm_config_db #(int)::set(null,"*","PORT_1635_COUNT",port_count[1635]);
       uvm_config_db #(int)::set(null,"*","PORT_1636_COUNT",port_count[1636]);
       uvm_config_db #(int)::set(null,"*","PORT_1637_COUNT",port_count[1637]);
       uvm_config_db #(int)::set(null,"*","PORT_1638_COUNT",port_count[1638]);
       uvm_config_db #(int)::set(null,"*","PORT_1639_COUNT",port_count[1639]);
       uvm_config_db #(int)::set(null,"*","PORT_1640_COUNT",port_count[1640]);
       uvm_config_db #(int)::set(null,"*","PORT_1641_COUNT",port_count[1641]);
       uvm_config_db #(int)::set(null,"*","PORT_1642_COUNT",port_count[1642]);
       uvm_config_db #(int)::set(null,"*","PORT_1643_COUNT",port_count[1643]);
       uvm_config_db #(int)::set(null,"*","PORT_1644_COUNT",port_count[1644]);
       uvm_config_db #(int)::set(null,"*","PORT_1645_COUNT",port_count[1645]);
       uvm_config_db #(int)::set(null,"*","PORT_1646_COUNT",port_count[1646]);
       uvm_config_db #(int)::set(null,"*","PORT_1647_COUNT",port_count[1647]);
       uvm_config_db #(int)::set(null,"*","PORT_1648_COUNT",port_count[1648]);
       uvm_config_db #(int)::set(null,"*","PORT_1649_COUNT",port_count[1649]);
       uvm_config_db #(int)::set(null,"*","PORT_1650_COUNT",port_count[1650]);
       uvm_config_db #(int)::set(null,"*","PORT_1651_COUNT",port_count[1651]);
       uvm_config_db #(int)::set(null,"*","PORT_1652_COUNT",port_count[1652]);
       uvm_config_db #(int)::set(null,"*","PORT_1653_COUNT",port_count[1653]);
       uvm_config_db #(int)::set(null,"*","PORT_1654_COUNT",port_count[1654]);
       uvm_config_db #(int)::set(null,"*","PORT_1655_COUNT",port_count[1655]);
       uvm_config_db #(int)::set(null,"*","PORT_1656_COUNT",port_count[1656]);
       uvm_config_db #(int)::set(null,"*","PORT_1657_COUNT",port_count[1657]);
       uvm_config_db #(int)::set(null,"*","PORT_1658_COUNT",port_count[1658]);
       uvm_config_db #(int)::set(null,"*","PORT_1659_COUNT",port_count[1659]);
       uvm_config_db #(int)::set(null,"*","PORT_1660_COUNT",port_count[1660]);
       uvm_config_db #(int)::set(null,"*","PORT_1661_COUNT",port_count[1661]);
       uvm_config_db #(int)::set(null,"*","PORT_1662_COUNT",port_count[1662]);
       uvm_config_db #(int)::set(null,"*","PORT_1663_COUNT",port_count[1663]);
       uvm_config_db #(int)::set(null,"*","PORT_1664_COUNT",port_count[1664]);
       uvm_config_db #(int)::set(null,"*","PORT_1665_COUNT",port_count[1665]);
       uvm_config_db #(int)::set(null,"*","PORT_1666_COUNT",port_count[1666]);
       uvm_config_db #(int)::set(null,"*","PORT_1667_COUNT",port_count[1667]);
       uvm_config_db #(int)::set(null,"*","PORT_1668_COUNT",port_count[1668]);
       uvm_config_db #(int)::set(null,"*","PORT_1669_COUNT",port_count[1669]);
       uvm_config_db #(int)::set(null,"*","PORT_1670_COUNT",port_count[1670]);
       uvm_config_db #(int)::set(null,"*","PORT_1671_COUNT",port_count[1671]);
       uvm_config_db #(int)::set(null,"*","PORT_1672_COUNT",port_count[1672]);
       uvm_config_db #(int)::set(null,"*","PORT_1673_COUNT",port_count[1673]);
       uvm_config_db #(int)::set(null,"*","PORT_1674_COUNT",port_count[1674]);
       uvm_config_db #(int)::set(null,"*","PORT_1675_COUNT",port_count[1675]);
       uvm_config_db #(int)::set(null,"*","PORT_1676_COUNT",port_count[1676]);
       uvm_config_db #(int)::set(null,"*","PORT_1677_COUNT",port_count[1677]);
       uvm_config_db #(int)::set(null,"*","PORT_1678_COUNT",port_count[1678]);
       uvm_config_db #(int)::set(null,"*","PORT_1679_COUNT",port_count[1679]);
       uvm_config_db #(int)::set(null,"*","PORT_1680_COUNT",port_count[1680]);
       uvm_config_db #(int)::set(null,"*","PORT_1681_COUNT",port_count[1681]);
       uvm_config_db #(int)::set(null,"*","PORT_1682_COUNT",port_count[1682]);
       uvm_config_db #(int)::set(null,"*","PORT_1683_COUNT",port_count[1683]);
       uvm_config_db #(int)::set(null,"*","PORT_1684_COUNT",port_count[1684]);
       uvm_config_db #(int)::set(null,"*","PORT_1685_COUNT",port_count[1685]);
       uvm_config_db #(int)::set(null,"*","PORT_1686_COUNT",port_count[1686]);
       uvm_config_db #(int)::set(null,"*","PORT_1687_COUNT",port_count[1687]);
       uvm_config_db #(int)::set(null,"*","PORT_1688_COUNT",port_count[1688]);
       uvm_config_db #(int)::set(null,"*","PORT_1689_COUNT",port_count[1689]);
       uvm_config_db #(int)::set(null,"*","PORT_1690_COUNT",port_count[1690]);
       uvm_config_db #(int)::set(null,"*","PORT_1691_COUNT",port_count[1691]);
       uvm_config_db #(int)::set(null,"*","PORT_1692_COUNT",port_count[1692]);
       uvm_config_db #(int)::set(null,"*","PORT_1693_COUNT",port_count[1693]);
       uvm_config_db #(int)::set(null,"*","PORT_1694_COUNT",port_count[1694]);
       uvm_config_db #(int)::set(null,"*","PORT_1695_COUNT",port_count[1695]);
       uvm_config_db #(int)::set(null,"*","PORT_1696_COUNT",port_count[1696]);
       uvm_config_db #(int)::set(null,"*","PORT_1697_COUNT",port_count[1697]);
       uvm_config_db #(int)::set(null,"*","PORT_1698_COUNT",port_count[1698]);
       uvm_config_db #(int)::set(null,"*","PORT_1699_COUNT",port_count[1699]);
       uvm_config_db #(int)::set(null,"*","PORT_1700_COUNT",port_count[1700]);
       uvm_config_db #(int)::set(null,"*","PORT_1701_COUNT",port_count[1701]);
       uvm_config_db #(int)::set(null,"*","PORT_1702_COUNT",port_count[1702]);
       uvm_config_db #(int)::set(null,"*","PORT_1703_COUNT",port_count[1703]);
       uvm_config_db #(int)::set(null,"*","PORT_1704_COUNT",port_count[1704]);
       uvm_config_db #(int)::set(null,"*","PORT_1705_COUNT",port_count[1705]);
       uvm_config_db #(int)::set(null,"*","PORT_1706_COUNT",port_count[1706]);
       uvm_config_db #(int)::set(null,"*","PORT_1707_COUNT",port_count[1707]);
       uvm_config_db #(int)::set(null,"*","PORT_1708_COUNT",port_count[1708]);
       uvm_config_db #(int)::set(null,"*","PORT_1709_COUNT",port_count[1709]);
       uvm_config_db #(int)::set(null,"*","PORT_1710_COUNT",port_count[1710]);
       uvm_config_db #(int)::set(null,"*","PORT_1711_COUNT",port_count[1711]);
       uvm_config_db #(int)::set(null,"*","PORT_1712_COUNT",port_count[1712]);
       uvm_config_db #(int)::set(null,"*","PORT_1713_COUNT",port_count[1713]);
       uvm_config_db #(int)::set(null,"*","PORT_1714_COUNT",port_count[1714]);
       uvm_config_db #(int)::set(null,"*","PORT_1715_COUNT",port_count[1715]);
       uvm_config_db #(int)::set(null,"*","PORT_1716_COUNT",port_count[1716]);
       uvm_config_db #(int)::set(null,"*","PORT_1717_COUNT",port_count[1717]);
       uvm_config_db #(int)::set(null,"*","PORT_1718_COUNT",port_count[1718]);
       uvm_config_db #(int)::set(null,"*","PORT_1719_COUNT",port_count[1719]);
       uvm_config_db #(int)::set(null,"*","PORT_1720_COUNT",port_count[1720]);
       uvm_config_db #(int)::set(null,"*","PORT_1721_COUNT",port_count[1721]);
       uvm_config_db #(int)::set(null,"*","PORT_1722_COUNT",port_count[1722]);
       uvm_config_db #(int)::set(null,"*","PORT_1723_COUNT",port_count[1723]);
       uvm_config_db #(int)::set(null,"*","PORT_1724_COUNT",port_count[1724]);
       uvm_config_db #(int)::set(null,"*","PORT_1725_COUNT",port_count[1725]);
       uvm_config_db #(int)::set(null,"*","PORT_1726_COUNT",port_count[1726]);
       uvm_config_db #(int)::set(null,"*","PORT_1727_COUNT",port_count[1727]);
       uvm_config_db #(int)::set(null,"*","PORT_1728_COUNT",port_count[1728]);
       uvm_config_db #(int)::set(null,"*","PORT_1729_COUNT",port_count[1729]);
       uvm_config_db #(int)::set(null,"*","PORT_1730_COUNT",port_count[1730]);
       uvm_config_db #(int)::set(null,"*","PORT_1731_COUNT",port_count[1731]);
       uvm_config_db #(int)::set(null,"*","PORT_1732_COUNT",port_count[1732]);
       uvm_config_db #(int)::set(null,"*","PORT_1733_COUNT",port_count[1733]);
       uvm_config_db #(int)::set(null,"*","PORT_1734_COUNT",port_count[1734]);
       uvm_config_db #(int)::set(null,"*","PORT_1735_COUNT",port_count[1735]);
       uvm_config_db #(int)::set(null,"*","PORT_1736_COUNT",port_count[1736]);
       uvm_config_db #(int)::set(null,"*","PORT_1737_COUNT",port_count[1737]);
       uvm_config_db #(int)::set(null,"*","PORT_1738_COUNT",port_count[1738]);
       uvm_config_db #(int)::set(null,"*","PORT_1739_COUNT",port_count[1739]);
       uvm_config_db #(int)::set(null,"*","PORT_1740_COUNT",port_count[1740]);
       uvm_config_db #(int)::set(null,"*","PORT_1741_COUNT",port_count[1741]);
       uvm_config_db #(int)::set(null,"*","PORT_1742_COUNT",port_count[1742]);
       uvm_config_db #(int)::set(null,"*","PORT_1743_COUNT",port_count[1743]);
       uvm_config_db #(int)::set(null,"*","PORT_1744_COUNT",port_count[1744]);
       uvm_config_db #(int)::set(null,"*","PORT_1745_COUNT",port_count[1745]);
       uvm_config_db #(int)::set(null,"*","PORT_1746_COUNT",port_count[1746]);
       uvm_config_db #(int)::set(null,"*","PORT_1747_COUNT",port_count[1747]);
       uvm_config_db #(int)::set(null,"*","PORT_1748_COUNT",port_count[1748]);
       uvm_config_db #(int)::set(null,"*","PORT_1749_COUNT",port_count[1749]);
       uvm_config_db #(int)::set(null,"*","PORT_1750_COUNT",port_count[1750]);
       uvm_config_db #(int)::set(null,"*","PORT_1751_COUNT",port_count[1751]);
       uvm_config_db #(int)::set(null,"*","PORT_1752_COUNT",port_count[1752]);
       uvm_config_db #(int)::set(null,"*","PORT_1753_COUNT",port_count[1753]);
       uvm_config_db #(int)::set(null,"*","PORT_1754_COUNT",port_count[1754]);
       uvm_config_db #(int)::set(null,"*","PORT_1755_COUNT",port_count[1755]);
       uvm_config_db #(int)::set(null,"*","PORT_1756_COUNT",port_count[1756]);
       uvm_config_db #(int)::set(null,"*","PORT_1757_COUNT",port_count[1757]);
       uvm_config_db #(int)::set(null,"*","PORT_1758_COUNT",port_count[1758]);
       uvm_config_db #(int)::set(null,"*","PORT_1759_COUNT",port_count[1759]);
       uvm_config_db #(int)::set(null,"*","PORT_1760_COUNT",port_count[1760]);
       uvm_config_db #(int)::set(null,"*","PORT_1761_COUNT",port_count[1761]);
       uvm_config_db #(int)::set(null,"*","PORT_1762_COUNT",port_count[1762]);
       uvm_config_db #(int)::set(null,"*","PORT_1763_COUNT",port_count[1763]);
       uvm_config_db #(int)::set(null,"*","PORT_1764_COUNT",port_count[1764]);
       uvm_config_db #(int)::set(null,"*","PORT_1765_COUNT",port_count[1765]);
       uvm_config_db #(int)::set(null,"*","PORT_1766_COUNT",port_count[1766]);
       uvm_config_db #(int)::set(null,"*","PORT_1767_COUNT",port_count[1767]);
       uvm_config_db #(int)::set(null,"*","PORT_1768_COUNT",port_count[1768]);
       uvm_config_db #(int)::set(null,"*","PORT_1769_COUNT",port_count[1769]);
       uvm_config_db #(int)::set(null,"*","PORT_1770_COUNT",port_count[1770]);
       uvm_config_db #(int)::set(null,"*","PORT_1771_COUNT",port_count[1771]);
       uvm_config_db #(int)::set(null,"*","PORT_1772_COUNT",port_count[1772]);
       uvm_config_db #(int)::set(null,"*","PORT_1773_COUNT",port_count[1773]);
       uvm_config_db #(int)::set(null,"*","PORT_1774_COUNT",port_count[1774]);
       uvm_config_db #(int)::set(null,"*","PORT_1775_COUNT",port_count[1775]);
       uvm_config_db #(int)::set(null,"*","PORT_1776_COUNT",port_count[1776]);
       uvm_config_db #(int)::set(null,"*","PORT_1777_COUNT",port_count[1777]);
       uvm_config_db #(int)::set(null,"*","PORT_1778_COUNT",port_count[1778]);
       uvm_config_db #(int)::set(null,"*","PORT_1779_COUNT",port_count[1779]);
       uvm_config_db #(int)::set(null,"*","PORT_1780_COUNT",port_count[1780]);
       uvm_config_db #(int)::set(null,"*","PORT_1781_COUNT",port_count[1781]);
       uvm_config_db #(int)::set(null,"*","PORT_1782_COUNT",port_count[1782]);
       uvm_config_db #(int)::set(null,"*","PORT_1783_COUNT",port_count[1783]);
       uvm_config_db #(int)::set(null,"*","PORT_1784_COUNT",port_count[1784]);
       uvm_config_db #(int)::set(null,"*","PORT_1785_COUNT",port_count[1785]);
       uvm_config_db #(int)::set(null,"*","PORT_1786_COUNT",port_count[1786]);
       uvm_config_db #(int)::set(null,"*","PORT_1787_COUNT",port_count[1787]);
       uvm_config_db #(int)::set(null,"*","PORT_1788_COUNT",port_count[1788]);
       uvm_config_db #(int)::set(null,"*","PORT_1789_COUNT",port_count[1789]);
       uvm_config_db #(int)::set(null,"*","PORT_1790_COUNT",port_count[1790]);
       uvm_config_db #(int)::set(null,"*","PORT_1791_COUNT",port_count[1791]);
       uvm_config_db #(int)::set(null,"*","PORT_1792_COUNT",port_count[1792]);
       uvm_config_db #(int)::set(null,"*","PORT_1793_COUNT",port_count[1793]);
       uvm_config_db #(int)::set(null,"*","PORT_1794_COUNT",port_count[1794]);
       uvm_config_db #(int)::set(null,"*","PORT_1795_COUNT",port_count[1795]);
       uvm_config_db #(int)::set(null,"*","PORT_1796_COUNT",port_count[1796]);
       uvm_config_db #(int)::set(null,"*","PORT_1797_COUNT",port_count[1797]);
       uvm_config_db #(int)::set(null,"*","PORT_1798_COUNT",port_count[1798]);
       uvm_config_db #(int)::set(null,"*","PORT_1799_COUNT",port_count[1799]);
       uvm_config_db #(int)::set(null,"*","PORT_1800_COUNT",port_count[1800]);
       uvm_config_db #(int)::set(null,"*","PORT_1801_COUNT",port_count[1801]);
       uvm_config_db #(int)::set(null,"*","PORT_1802_COUNT",port_count[1802]);
       uvm_config_db #(int)::set(null,"*","PORT_1803_COUNT",port_count[1803]);
       uvm_config_db #(int)::set(null,"*","PORT_1804_COUNT",port_count[1804]);
       uvm_config_db #(int)::set(null,"*","PORT_1805_COUNT",port_count[1805]);
       uvm_config_db #(int)::set(null,"*","PORT_1806_COUNT",port_count[1806]);
       uvm_config_db #(int)::set(null,"*","PORT_1807_COUNT",port_count[1807]);
       uvm_config_db #(int)::set(null,"*","PORT_1808_COUNT",port_count[1808]);
       uvm_config_db #(int)::set(null,"*","PORT_1809_COUNT",port_count[1809]);
       uvm_config_db #(int)::set(null,"*","PORT_1810_COUNT",port_count[1810]);
       uvm_config_db #(int)::set(null,"*","PORT_1811_COUNT",port_count[1811]);
       uvm_config_db #(int)::set(null,"*","PORT_1812_COUNT",port_count[1812]);
       uvm_config_db #(int)::set(null,"*","PORT_1813_COUNT",port_count[1813]);
       uvm_config_db #(int)::set(null,"*","PORT_1814_COUNT",port_count[1814]);
       uvm_config_db #(int)::set(null,"*","PORT_1815_COUNT",port_count[1815]);
       uvm_config_db #(int)::set(null,"*","PORT_1816_COUNT",port_count[1816]);
       uvm_config_db #(int)::set(null,"*","PORT_1817_COUNT",port_count[1817]);
       uvm_config_db #(int)::set(null,"*","PORT_1818_COUNT",port_count[1818]);
       uvm_config_db #(int)::set(null,"*","PORT_1819_COUNT",port_count[1819]);
       uvm_config_db #(int)::set(null,"*","PORT_1820_COUNT",port_count[1820]);
       uvm_config_db #(int)::set(null,"*","PORT_1821_COUNT",port_count[1821]);
       uvm_config_db #(int)::set(null,"*","PORT_1822_COUNT",port_count[1822]);
       uvm_config_db #(int)::set(null,"*","PORT_1823_COUNT",port_count[1823]);
       uvm_config_db #(int)::set(null,"*","PORT_1824_COUNT",port_count[1824]);
       uvm_config_db #(int)::set(null,"*","PORT_1825_COUNT",port_count[1825]);
       uvm_config_db #(int)::set(null,"*","PORT_1826_COUNT",port_count[1826]);
       uvm_config_db #(int)::set(null,"*","PORT_1827_COUNT",port_count[1827]);
       uvm_config_db #(int)::set(null,"*","PORT_1828_COUNT",port_count[1828]);
       uvm_config_db #(int)::set(null,"*","PORT_1829_COUNT",port_count[1829]);
       uvm_config_db #(int)::set(null,"*","PORT_1830_COUNT",port_count[1830]);
       uvm_config_db #(int)::set(null,"*","PORT_1831_COUNT",port_count[1831]);
       uvm_config_db #(int)::set(null,"*","PORT_1832_COUNT",port_count[1832]);
       uvm_config_db #(int)::set(null,"*","PORT_1833_COUNT",port_count[1833]);
       uvm_config_db #(int)::set(null,"*","PORT_1834_COUNT",port_count[1834]);
       uvm_config_db #(int)::set(null,"*","PORT_1835_COUNT",port_count[1835]);
       uvm_config_db #(int)::set(null,"*","PORT_1836_COUNT",port_count[1836]);
       uvm_config_db #(int)::set(null,"*","PORT_1837_COUNT",port_count[1837]);
       uvm_config_db #(int)::set(null,"*","PORT_1838_COUNT",port_count[1838]);
       uvm_config_db #(int)::set(null,"*","PORT_1839_COUNT",port_count[1839]);
       uvm_config_db #(int)::set(null,"*","PORT_1840_COUNT",port_count[1840]);
       uvm_config_db #(int)::set(null,"*","PORT_1841_COUNT",port_count[1841]);
       uvm_config_db #(int)::set(null,"*","PORT_1842_COUNT",port_count[1842]);
       uvm_config_db #(int)::set(null,"*","PORT_1843_COUNT",port_count[1843]);
       uvm_config_db #(int)::set(null,"*","PORT_1844_COUNT",port_count[1844]);
       uvm_config_db #(int)::set(null,"*","PORT_1845_COUNT",port_count[1845]);
       uvm_config_db #(int)::set(null,"*","PORT_1846_COUNT",port_count[1846]);
       uvm_config_db #(int)::set(null,"*","PORT_1847_COUNT",port_count[1847]);
       uvm_config_db #(int)::set(null,"*","PORT_1848_COUNT",port_count[1848]);
       uvm_config_db #(int)::set(null,"*","PORT_1849_COUNT",port_count[1849]);
       uvm_config_db #(int)::set(null,"*","PORT_1850_COUNT",port_count[1850]);
       uvm_config_db #(int)::set(null,"*","PORT_1851_COUNT",port_count[1851]);
       uvm_config_db #(int)::set(null,"*","PORT_1852_COUNT",port_count[1852]);
       uvm_config_db #(int)::set(null,"*","PORT_1853_COUNT",port_count[1853]);
       uvm_config_db #(int)::set(null,"*","PORT_1854_COUNT",port_count[1854]);
       uvm_config_db #(int)::set(null,"*","PORT_1855_COUNT",port_count[1855]);
       uvm_config_db #(int)::set(null,"*","PORT_1856_COUNT",port_count[1856]);
       uvm_config_db #(int)::set(null,"*","PORT_1857_COUNT",port_count[1857]);
       uvm_config_db #(int)::set(null,"*","PORT_1858_COUNT",port_count[1858]);
       uvm_config_db #(int)::set(null,"*","PORT_1859_COUNT",port_count[1859]);
       uvm_config_db #(int)::set(null,"*","PORT_1860_COUNT",port_count[1860]);
       uvm_config_db #(int)::set(null,"*","PORT_1861_COUNT",port_count[1861]);
       uvm_config_db #(int)::set(null,"*","PORT_1862_COUNT",port_count[1862]);
       uvm_config_db #(int)::set(null,"*","PORT_1863_COUNT",port_count[1863]);
       uvm_config_db #(int)::set(null,"*","PORT_1864_COUNT",port_count[1864]);
       uvm_config_db #(int)::set(null,"*","PORT_1865_COUNT",port_count[1865]);
       uvm_config_db #(int)::set(null,"*","PORT_1866_COUNT",port_count[1866]);
       uvm_config_db #(int)::set(null,"*","PORT_1867_COUNT",port_count[1867]);
       uvm_config_db #(int)::set(null,"*","PORT_1868_COUNT",port_count[1868]);
       uvm_config_db #(int)::set(null,"*","PORT_1869_COUNT",port_count[1869]);
       uvm_config_db #(int)::set(null,"*","PORT_1870_COUNT",port_count[1870]);
       uvm_config_db #(int)::set(null,"*","PORT_1871_COUNT",port_count[1871]);
       uvm_config_db #(int)::set(null,"*","PORT_1872_COUNT",port_count[1872]);
       uvm_config_db #(int)::set(null,"*","PORT_1873_COUNT",port_count[1873]);
       uvm_config_db #(int)::set(null,"*","PORT_1874_COUNT",port_count[1874]);
       uvm_config_db #(int)::set(null,"*","PORT_1875_COUNT",port_count[1875]);
       uvm_config_db #(int)::set(null,"*","PORT_1876_COUNT",port_count[1876]);
       uvm_config_db #(int)::set(null,"*","PORT_1877_COUNT",port_count[1877]);
       uvm_config_db #(int)::set(null,"*","PORT_1878_COUNT",port_count[1878]);
       uvm_config_db #(int)::set(null,"*","PORT_1879_COUNT",port_count[1879]);
       uvm_config_db #(int)::set(null,"*","PORT_1880_COUNT",port_count[1880]);
       uvm_config_db #(int)::set(null,"*","PORT_1881_COUNT",port_count[1881]);
       uvm_config_db #(int)::set(null,"*","PORT_1882_COUNT",port_count[1882]);
       uvm_config_db #(int)::set(null,"*","PORT_1883_COUNT",port_count[1883]);
       uvm_config_db #(int)::set(null,"*","PORT_1884_COUNT",port_count[1884]);
       uvm_config_db #(int)::set(null,"*","PORT_1885_COUNT",port_count[1885]);
       uvm_config_db #(int)::set(null,"*","PORT_1886_COUNT",port_count[1886]);
       uvm_config_db #(int)::set(null,"*","PORT_1887_COUNT",port_count[1887]);
       uvm_config_db #(int)::set(null,"*","PORT_1888_COUNT",port_count[1888]);
       uvm_config_db #(int)::set(null,"*","PORT_1889_COUNT",port_count[1889]);
       uvm_config_db #(int)::set(null,"*","PORT_1890_COUNT",port_count[1890]);
       uvm_config_db #(int)::set(null,"*","PORT_1891_COUNT",port_count[1891]);
       uvm_config_db #(int)::set(null,"*","PORT_1892_COUNT",port_count[1892]);
       uvm_config_db #(int)::set(null,"*","PORT_1893_COUNT",port_count[1893]);
       uvm_config_db #(int)::set(null,"*","PORT_1894_COUNT",port_count[1894]);
       uvm_config_db #(int)::set(null,"*","PORT_1895_COUNT",port_count[1895]);
       uvm_config_db #(int)::set(null,"*","PORT_1896_COUNT",port_count[1896]);
       uvm_config_db #(int)::set(null,"*","PORT_1897_COUNT",port_count[1897]);
       uvm_config_db #(int)::set(null,"*","PORT_1898_COUNT",port_count[1898]);
       uvm_config_db #(int)::set(null,"*","PORT_1899_COUNT",port_count[1899]);
       uvm_config_db #(int)::set(null,"*","PORT_1900_COUNT",port_count[1900]);
       uvm_config_db #(int)::set(null,"*","PORT_1901_COUNT",port_count[1901]);
       uvm_config_db #(int)::set(null,"*","PORT_1902_COUNT",port_count[1902]);
       uvm_config_db #(int)::set(null,"*","PORT_1903_COUNT",port_count[1903]);
       uvm_config_db #(int)::set(null,"*","PORT_1904_COUNT",port_count[1904]);
       uvm_config_db #(int)::set(null,"*","PORT_1905_COUNT",port_count[1905]);
       uvm_config_db #(int)::set(null,"*","PORT_1906_COUNT",port_count[1906]);
       uvm_config_db #(int)::set(null,"*","PORT_1907_COUNT",port_count[1907]);
       uvm_config_db #(int)::set(null,"*","PORT_1908_COUNT",port_count[1908]);
       uvm_config_db #(int)::set(null,"*","PORT_1909_COUNT",port_count[1909]);
       uvm_config_db #(int)::set(null,"*","PORT_1910_COUNT",port_count[1910]);
       uvm_config_db #(int)::set(null,"*","PORT_1911_COUNT",port_count[1911]);
       uvm_config_db #(int)::set(null,"*","PORT_1912_COUNT",port_count[1912]);
       uvm_config_db #(int)::set(null,"*","PORT_1913_COUNT",port_count[1913]);
       uvm_config_db #(int)::set(null,"*","PORT_1914_COUNT",port_count[1914]);
       uvm_config_db #(int)::set(null,"*","PORT_1915_COUNT",port_count[1915]);
       uvm_config_db #(int)::set(null,"*","PORT_1916_COUNT",port_count[1916]);
       uvm_config_db #(int)::set(null,"*","PORT_1917_COUNT",port_count[1917]);
       uvm_config_db #(int)::set(null,"*","PORT_1918_COUNT",port_count[1918]);
       uvm_config_db #(int)::set(null,"*","PORT_1919_COUNT",port_count[1919]);
       uvm_config_db #(int)::set(null,"*","PORT_1920_COUNT",port_count[1920]);
       uvm_config_db #(int)::set(null,"*","PORT_1921_COUNT",port_count[1921]);
       uvm_config_db #(int)::set(null,"*","PORT_1922_COUNT",port_count[1922]);
       uvm_config_db #(int)::set(null,"*","PORT_1923_COUNT",port_count[1923]);
       uvm_config_db #(int)::set(null,"*","PORT_1924_COUNT",port_count[1924]);
       uvm_config_db #(int)::set(null,"*","PORT_1925_COUNT",port_count[1925]);
       uvm_config_db #(int)::set(null,"*","PORT_1926_COUNT",port_count[1926]);
       uvm_config_db #(int)::set(null,"*","PORT_1927_COUNT",port_count[1927]);
       uvm_config_db #(int)::set(null,"*","PORT_1928_COUNT",port_count[1928]);
       uvm_config_db #(int)::set(null,"*","PORT_1929_COUNT",port_count[1929]);
       uvm_config_db #(int)::set(null,"*","PORT_1930_COUNT",port_count[1930]);
       uvm_config_db #(int)::set(null,"*","PORT_1931_COUNT",port_count[1931]);
       uvm_config_db #(int)::set(null,"*","PORT_1932_COUNT",port_count[1932]);
       uvm_config_db #(int)::set(null,"*","PORT_1933_COUNT",port_count[1933]);
       uvm_config_db #(int)::set(null,"*","PORT_1934_COUNT",port_count[1934]);
       uvm_config_db #(int)::set(null,"*","PORT_1935_COUNT",port_count[1935]);
       uvm_config_db #(int)::set(null,"*","PORT_1936_COUNT",port_count[1936]);
       uvm_config_db #(int)::set(null,"*","PORT_1937_COUNT",port_count[1937]);
       uvm_config_db #(int)::set(null,"*","PORT_1938_COUNT",port_count[1938]);
       uvm_config_db #(int)::set(null,"*","PORT_1939_COUNT",port_count[1939]);
       uvm_config_db #(int)::set(null,"*","PORT_1940_COUNT",port_count[1940]);
       uvm_config_db #(int)::set(null,"*","PORT_1941_COUNT",port_count[1941]);
       uvm_config_db #(int)::set(null,"*","PORT_1942_COUNT",port_count[1942]);
       uvm_config_db #(int)::set(null,"*","PORT_1943_COUNT",port_count[1943]);
       uvm_config_db #(int)::set(null,"*","PORT_1944_COUNT",port_count[1944]);
       uvm_config_db #(int)::set(null,"*","PORT_1945_COUNT",port_count[1945]);
       uvm_config_db #(int)::set(null,"*","PORT_1946_COUNT",port_count[1946]);
       uvm_config_db #(int)::set(null,"*","PORT_1947_COUNT",port_count[1947]);
       uvm_config_db #(int)::set(null,"*","PORT_1948_COUNT",port_count[1948]);
       uvm_config_db #(int)::set(null,"*","PORT_1949_COUNT",port_count[1949]);
       uvm_config_db #(int)::set(null,"*","PORT_1950_COUNT",port_count[1950]);
       uvm_config_db #(int)::set(null,"*","PORT_1951_COUNT",port_count[1951]);
       uvm_config_db #(int)::set(null,"*","PORT_1952_COUNT",port_count[1952]);
       uvm_config_db #(int)::set(null,"*","PORT_1953_COUNT",port_count[1953]);
       uvm_config_db #(int)::set(null,"*","PORT_1954_COUNT",port_count[1954]);
       uvm_config_db #(int)::set(null,"*","PORT_1955_COUNT",port_count[1955]);
       uvm_config_db #(int)::set(null,"*","PORT_1956_COUNT",port_count[1956]);
       uvm_config_db #(int)::set(null,"*","PORT_1957_COUNT",port_count[1957]);
       uvm_config_db #(int)::set(null,"*","PORT_1958_COUNT",port_count[1958]);
       uvm_config_db #(int)::set(null,"*","PORT_1959_COUNT",port_count[1959]);
       uvm_config_db #(int)::set(null,"*","PORT_1960_COUNT",port_count[1960]);
       uvm_config_db #(int)::set(null,"*","PORT_1961_COUNT",port_count[1961]);
       uvm_config_db #(int)::set(null,"*","PORT_1962_COUNT",port_count[1962]);
       uvm_config_db #(int)::set(null,"*","PORT_1963_COUNT",port_count[1963]);
       uvm_config_db #(int)::set(null,"*","PORT_1964_COUNT",port_count[1964]);
       uvm_config_db #(int)::set(null,"*","PORT_1965_COUNT",port_count[1965]);
       uvm_config_db #(int)::set(null,"*","PORT_1966_COUNT",port_count[1966]);
       uvm_config_db #(int)::set(null,"*","PORT_1967_COUNT",port_count[1967]);
       uvm_config_db #(int)::set(null,"*","PORT_1968_COUNT",port_count[1968]);
       uvm_config_db #(int)::set(null,"*","PORT_1969_COUNT",port_count[1969]);
       uvm_config_db #(int)::set(null,"*","PORT_1970_COUNT",port_count[1970]);
       uvm_config_db #(int)::set(null,"*","PORT_1971_COUNT",port_count[1971]);
       uvm_config_db #(int)::set(null,"*","PORT_1972_COUNT",port_count[1972]);
       uvm_config_db #(int)::set(null,"*","PORT_1973_COUNT",port_count[1973]);
       uvm_config_db #(int)::set(null,"*","PORT_1974_COUNT",port_count[1974]);
       uvm_config_db #(int)::set(null,"*","PORT_1975_COUNT",port_count[1975]);
       uvm_config_db #(int)::set(null,"*","PORT_1976_COUNT",port_count[1976]);
       uvm_config_db #(int)::set(null,"*","PORT_1977_COUNT",port_count[1977]);
       uvm_config_db #(int)::set(null,"*","PORT_1978_COUNT",port_count[1978]);
       uvm_config_db #(int)::set(null,"*","PORT_1979_COUNT",port_count[1979]);
       uvm_config_db #(int)::set(null,"*","PORT_1980_COUNT",port_count[1980]);
       uvm_config_db #(int)::set(null,"*","PORT_1981_COUNT",port_count[1981]);
       uvm_config_db #(int)::set(null,"*","PORT_1982_COUNT",port_count[1982]);
       uvm_config_db #(int)::set(null,"*","PORT_1983_COUNT",port_count[1983]);
       uvm_config_db #(int)::set(null,"*","PORT_1984_COUNT",port_count[1984]);
       uvm_config_db #(int)::set(null,"*","PORT_1985_COUNT",port_count[1985]);
       uvm_config_db #(int)::set(null,"*","PORT_1986_COUNT",port_count[1986]);
       uvm_config_db #(int)::set(null,"*","PORT_1987_COUNT",port_count[1987]);
       uvm_config_db #(int)::set(null,"*","PORT_1988_COUNT",port_count[1988]);
       uvm_config_db #(int)::set(null,"*","PORT_1989_COUNT",port_count[1989]);
       uvm_config_db #(int)::set(null,"*","PORT_1990_COUNT",port_count[1990]);
       uvm_config_db #(int)::set(null,"*","PORT_1991_COUNT",port_count[1991]);
       uvm_config_db #(int)::set(null,"*","PORT_1992_COUNT",port_count[1992]);
       uvm_config_db #(int)::set(null,"*","PORT_1993_COUNT",port_count[1993]);
       uvm_config_db #(int)::set(null,"*","PORT_1994_COUNT",port_count[1994]);
       uvm_config_db #(int)::set(null,"*","PORT_1995_COUNT",port_count[1995]);
       uvm_config_db #(int)::set(null,"*","PORT_1996_COUNT",port_count[1996]);
       uvm_config_db #(int)::set(null,"*","PORT_1997_COUNT",port_count[1997]);
       uvm_config_db #(int)::set(null,"*","PORT_1998_COUNT",port_count[1998]);
       uvm_config_db #(int)::set(null,"*","PORT_1999_COUNT",port_count[1999]);
       uvm_config_db #(int)::set(null,"*","PORT_2000_COUNT",port_count[2000]);
       uvm_config_db #(int)::set(null,"*","PORT_2001_COUNT",port_count[2001]);
       uvm_config_db #(int)::set(null,"*","PORT_2002_COUNT",port_count[2002]);
       uvm_config_db #(int)::set(null,"*","PORT_2003_COUNT",port_count[2003]);
       uvm_config_db #(int)::set(null,"*","PORT_2004_COUNT",port_count[2004]);
       uvm_config_db #(int)::set(null,"*","PORT_2005_COUNT",port_count[2005]);
       uvm_config_db #(int)::set(null,"*","PORT_2006_COUNT",port_count[2006]);
       uvm_config_db #(int)::set(null,"*","PORT_2007_COUNT",port_count[2007]);
       uvm_config_db #(int)::set(null,"*","PORT_2008_COUNT",port_count[2008]);
       uvm_config_db #(int)::set(null,"*","PORT_2009_COUNT",port_count[2009]);
       uvm_config_db #(int)::set(null,"*","PORT_2010_COUNT",port_count[2010]);
       uvm_config_db #(int)::set(null,"*","PORT_2011_COUNT",port_count[2011]);
       uvm_config_db #(int)::set(null,"*","PORT_2012_COUNT",port_count[2012]);
       uvm_config_db #(int)::set(null,"*","PORT_2013_COUNT",port_count[2013]);
       uvm_config_db #(int)::set(null,"*","PORT_2014_COUNT",port_count[2014]);
       uvm_config_db #(int)::set(null,"*","PORT_2015_COUNT",port_count[2015]);
       uvm_config_db #(int)::set(null,"*","PORT_2016_COUNT",port_count[2016]);
       uvm_config_db #(int)::set(null,"*","PORT_2017_COUNT",port_count[2017]);
       uvm_config_db #(int)::set(null,"*","PORT_2018_COUNT",port_count[2018]);
       uvm_config_db #(int)::set(null,"*","PORT_2019_COUNT",port_count[2019]);
       uvm_config_db #(int)::set(null,"*","PORT_2020_COUNT",port_count[2020]);
       uvm_config_db #(int)::set(null,"*","PORT_2021_COUNT",port_count[2021]);
       uvm_config_db #(int)::set(null,"*","PORT_2022_COUNT",port_count[2022]);
       uvm_config_db #(int)::set(null,"*","PORT_2023_COUNT",port_count[2023]);
       uvm_config_db #(int)::set(null,"*","PORT_2024_COUNT",port_count[2024]);
       uvm_config_db #(int)::set(null,"*","PORT_2025_COUNT",port_count[2025]);
       uvm_config_db #(int)::set(null,"*","PORT_2026_COUNT",port_count[2026]);
       uvm_config_db #(int)::set(null,"*","PORT_2027_COUNT",port_count[2027]);
       uvm_config_db #(int)::set(null,"*","PORT_2028_COUNT",port_count[2028]);
       uvm_config_db #(int)::set(null,"*","PORT_2029_COUNT",port_count[2029]);
       uvm_config_db #(int)::set(null,"*","PORT_2030_COUNT",port_count[2030]);
       uvm_config_db #(int)::set(null,"*","PORT_2031_COUNT",port_count[2031]);
       uvm_config_db #(int)::set(null,"*","PORT_2032_COUNT",port_count[2032]);
       uvm_config_db #(int)::set(null,"*","PORT_2033_COUNT",port_count[2033]);
       uvm_config_db #(int)::set(null,"*","PORT_2034_COUNT",port_count[2034]);
       uvm_config_db #(int)::set(null,"*","PORT_2035_COUNT",port_count[2035]);
       uvm_config_db #(int)::set(null,"*","PORT_2036_COUNT",port_count[2036]);
       uvm_config_db #(int)::set(null,"*","PORT_2037_COUNT",port_count[2037]);
       uvm_config_db #(int)::set(null,"*","PORT_2038_COUNT",port_count[2038]);
       uvm_config_db #(int)::set(null,"*","PORT_2039_COUNT",port_count[2039]);
       uvm_config_db #(int)::set(null,"*","PORT_2040_COUNT",port_count[2040]);
       uvm_config_db #(int)::set(null,"*","PORT_2041_COUNT",port_count[2041]);
       uvm_config_db #(int)::set(null,"*","PORT_2042_COUNT",port_count[2042]);
       uvm_config_db #(int)::set(null,"*","PORT_2043_COUNT",port_count[2043]);
       uvm_config_db #(int)::set(null,"*","PORT_2044_COUNT",port_count[2044]);
       uvm_config_db #(int)::set(null,"*","PORT_2045_COUNT",port_count[2045]);
       uvm_config_db #(int)::set(null,"*","PORT_2046_COUNT",port_count[2046]);
       uvm_config_db #(int)::set(null,"*","PORT_2047_COUNT",port_count[2047]);
       `endif

       `uvm_info(get_name(), "Exiting sequence...", UVM_LOW)
    endtask : body

endclass
