// Copyright (C) 2023 Intel Corporation
// SPDX-License-Identifier: MIT

`define TOP top_tb.pf_vf_mux_a

`define device_slave_connections(PORT) \
 force axis_if_D.slave_if[``PORT``].tvalid    =  `TOP.mx2fn_rx_port[``PORT``].tvalid        ;\
 force axis_if_D.slave_if[``PORT``].tlast     =  `TOP.mx2fn_rx_port[``PORT``].tlast         ;\
 force axis_if_D.slave_if[``PORT``].tuser     =  `TOP.mx2fn_rx_port[``PORT``].tuser_vendor  ;\
 force axis_if_D.slave_if[``PORT``].tdata     =  `TOP.mx2fn_rx_port[``PORT``].tdata         ;\
 force axis_if_D.slave_if[``PORT``].tkeep     =  `TOP.mx2fn_rx_port[``PORT``].tkeep         ;\
 force axis_if_D.slave_if[``PORT``].tready    =  `TOP.mx2fn_rx_port[``PORT``].tready        ;\
 force axis_if_D.slave_if[``PORT``].tready    =  1'b1        ;\
 force `TOP.fn2mx_tx_port[``PORT``].tvalid          =    axis_if_D.master_if[``PORT``].tvalid   ;\ 
 force `TOP.fn2mx_tx_port[``PORT``].tlast           =    axis_if_D.master_if[``PORT``].tlast    ;\   
 force `TOP.fn2mx_tx_port[``PORT``].tuser_vendor    =    axis_if_D.master_if[``PORT``].tuser    ;\   
 force `TOP.fn2mx_tx_port[``PORT``].tdata           =    axis_if_D.master_if[``PORT``].tdata    ;\   
 force `TOP.fn2mx_tx_port[``PORT``].tkeep           =    axis_if_D.master_if[``PORT``].tkeep    ;\   
 force axis_if_D.master_if[``PORT``].tready         =    `TOP.fn2mx_tx_port[``PORT``].tready    ;\


 `define device_slave_connections_N(RTL_PORT,VIP_PORT) \
 force axis_if_DN.slave_if[``VIP_PORT``].tvalid    =  `TOP.mx2fn_rx_port[``RTL_PORT``].tvalid        ;\
 force axis_if_DN.slave_if[``VIP_PORT``].tlast     =  `TOP.mx2fn_rx_port[``RTL_PORT``].tlast         ;\
 force axis_if_DN.slave_if[``VIP_PORT``].tuser     =  `TOP.mx2fn_rx_port[``RTL_PORT``].tuser_vendor  ;\
 force axis_if_DN.slave_if[``VIP_PORT``].tdata     =  `TOP.mx2fn_rx_port[``RTL_PORT``].tdata         ;\
 force axis_if_DN.slave_if[``VIP_PORT``].tkeep     =  `TOP.mx2fn_rx_port[``RTL_PORT``].tkeep         ;\
 force axis_if_DN.slave_if[``VIP_PORT``].tready    =  `TOP.mx2fn_rx_port[``RTL_PORT``].tready        ;\
 force axis_if_DN.slave_if[``VIP_PORT``].tready    =  1'b1        ;\
 force `TOP.fn2mx_tx_port[``RTL_PORT``].tvalid          =    axis_if_DN.master_if[``VIP_PORT``].tvalid   ;\ 
 force `TOP.fn2mx_tx_port[``RTL_PORT``].tlast           =    axis_if_DN.master_if[``VIP_PORT``].tlast    ;\   
 force `TOP.fn2mx_tx_port[``RTL_PORT``].tuser_vendor    =    axis_if_DN.master_if[``VIP_PORT``].tuser    ;\   
 force `TOP.fn2mx_tx_port[``RTL_PORT``].tdata           =    axis_if_DN.master_if[``VIP_PORT``].tdata    ;\   
 force `TOP.fn2mx_tx_port[``RTL_PORT``].tkeep           =    axis_if_DN.master_if[``VIP_PORT``].tkeep    ;\   
 force axis_if_DN.master_if[``VIP_PORT``].tready         =    `TOP.fn2mx_tx_port[``RTL_PORT``].tready    ;\

 `define device_slave_connections_TB_CONFIG_4(VIP_NUM,RTL_PORT,VIP_PORT) \
 force TB4_axis_if_D``VIP_NUM``.slave_if[``VIP_PORT``].tvalid    =  `TOP.mx2fn_rx_port[``RTL_PORT``].tvalid        ;\
 force TB4_axis_if_D``VIP_NUM``.slave_if[``VIP_PORT``].tlast     =  `TOP.mx2fn_rx_port[``RTL_PORT``].tlast         ;\
 force TB4_axis_if_D``VIP_NUM``.slave_if[``VIP_PORT``].tuser     =  `TOP.mx2fn_rx_port[``RTL_PORT``].tuser_vendor  ;\
 force TB4_axis_if_D``VIP_NUM``.slave_if[``VIP_PORT``].tdata     =  `TOP.mx2fn_rx_port[``RTL_PORT``].tdata         ;\
 force TB4_axis_if_D``VIP_NUM``.slave_if[``VIP_PORT``].tkeep     =  `TOP.mx2fn_rx_port[``RTL_PORT``].tkeep         ;\
 force TB4_axis_if_D``VIP_NUM``.slave_if[``VIP_PORT``].tready    =  `TOP.mx2fn_rx_port[``RTL_PORT``].tready        ;\
 force TB4_axis_if_D``VIP_NUM``.slave_if[``VIP_PORT``].tready    =  1'b1        ;\
 force `TOP.fn2mx_tx_port[``RTL_PORT``].tvalid          =    TB4_axis_if_D``VIP_NUM``.master_if[``VIP_PORT``].tvalid   ;\ 
 force `TOP.fn2mx_tx_port[``RTL_PORT``].tlast           =    TB4_axis_if_D``VIP_NUM``.master_if[``VIP_PORT``].tlast    ;\   
 force `TOP.fn2mx_tx_port[``RTL_PORT``].tuser_vendor    =    TB4_axis_if_D``VIP_NUM``.master_if[``VIP_PORT``].tuser    ;\   
 force `TOP.fn2mx_tx_port[``RTL_PORT``].tdata           =    TB4_axis_if_D``VIP_NUM``.master_if[``VIP_PORT``].tdata    ;\   
 force `TOP.fn2mx_tx_port[``RTL_PORT``].tkeep           =    TB4_axis_if_D``VIP_NUM``.master_if[``VIP_PORT``].tkeep    ;\   
 force TB4_axis_if_D``VIP_NUM``.master_if[``VIP_PORT``].tready         =    `TOP.fn2mx_tx_port[``RTL_PORT``].tready    ;\



`include "uvm_pkg.sv"
`ifdef TB_CONFIG_1
module AXI_VIP (svt_axi_if axis_if_D,axis_if_H);
`elsif TB_CONFIG_4
module AXI_VIP (svt_axi_if axis_if_D,axis_if_H,TB4_axis_if_D0,TB4_axis_if_D1,TB4_axis_if_D2,TB4_axis_if_D3);
`else
module AXI_VIP (svt_axi_if axis_if_D,axis_if_DN,axis_if_H);
`endif

import uvm_pkg::*;
bit      VA ; 
bit[3:0] VF ;
bit[2:0] PF ;
genvar i;

assign axis_if_H.common_aclk = `TOP.clk;
assign axis_if_H.master_if[0].aresetn = `TOP.rst_n;
assign axis_if_H.slave_if[0].aresetn = `TOP.rst_n; 

assign axis_if_D.common_aclk = `TOP.clk;
`ifndef TB_CONFIG_4
   for(i=0;i<16;i++) begin
     assign axis_if_D.slave_if[i].aresetn = `TOP.rst_n; 
     assign axis_if_D.master_if[i].aresetn = `TOP.rst_n;
   end  
`endif

`ifndef TB_CONFIG_1
  `ifdef TB_CONFIG_4
     assign TB4_axis_if_D0.common_aclk = `TOP.clk;
     assign TB4_axis_if_D1.common_aclk = `TOP.clk;
     assign TB4_axis_if_D2.common_aclk = `TOP.clk;
     assign TB4_axis_if_D3.common_aclk = `TOP.clk;
     for(i=0;i<450;i++) begin
        assign axis_if_D.slave_if[i].aresetn = `TOP.rst_n; 
        assign axis_if_D.master_if[i].aresetn = `TOP.rst_n;
        assign TB4_axis_if_D0.slave_if[i].aresetn = `TOP.rst_n; 
        assign TB4_axis_if_D0.master_if[i].aresetn = `TOP.rst_n;
        assign TB4_axis_if_D1.slave_if[i].aresetn = `TOP.rst_n; 
        assign TB4_axis_if_D1.master_if[i].aresetn = `TOP.rst_n;
        assign TB4_axis_if_D2.slave_if[i].aresetn = `TOP.rst_n; 
        assign TB4_axis_if_D2.master_if[i].aresetn = `TOP.rst_n;
        assign TB4_axis_if_D3.slave_if[i].aresetn = `TOP.rst_n; 
        assign TB4_axis_if_D3.master_if[i].aresetn = `TOP.rst_n;
     end
  `else
     assign axis_if_DN.common_aclk = `TOP.clk;
     for(i=0;i<16;i++) begin
       assign axis_if_DN.slave_if[i].aresetn = `TOP.rst_n; 
       assign axis_if_DN.master_if[i].aresetn = `TOP.rst_n;
     end
   `endif 
`endif

initial begin 

  //=======================
  // Host --> MUX 
  //=======================
  force `TOP.ho2mx_rx_port.tvalid         =  axis_if_H.master_if[0].tvalid;
  force `TOP.ho2mx_rx_port.tlast          =  axis_if_H.master_if[0].tlast;
  force `TOP.ho2mx_rx_port.tuser_vendor   =  axis_if_H.master_if[0].tuser;
  force `TOP.ho2mx_rx_port.tdata          =  axis_if_H.master_if[0].tdata;
  force `TOP.ho2mx_rx_port.tkeep          =  axis_if_H.master_if[0].tkeep;
  force axis_if_H.master_if[0].tready     = `TOP.ho2mx_rx_port.tready ; 

  //==============================================
  // Mux --> Device Slave and Device Master to Mux 
  //==============================================

  `device_slave_connections(0);
  `device_slave_connections(1);
  `device_slave_connections(2);
  `device_slave_connections(3);
  `device_slave_connections(4);
  `device_slave_connections(5);
  `device_slave_connections(6);
  `device_slave_connections(7);
  `device_slave_connections(8);
  `device_slave_connections(9);
  `device_slave_connections(10);
  `device_slave_connections(11);
  `device_slave_connections(12);
  `device_slave_connections(13);
  `device_slave_connections(14);
  `device_slave_connections(15);
 `ifdef TB_CONFIG_4
  `device_slave_connections(16);
  `device_slave_connections(17);
  `device_slave_connections(18);
  `device_slave_connections(19);
  `device_slave_connections(20);
  `device_slave_connections(21);
  `device_slave_connections(22);
  `device_slave_connections(23);
  `device_slave_connections(24);
  `device_slave_connections(25);
  `device_slave_connections(26);
  `device_slave_connections(27);
  `device_slave_connections(28);
  `device_slave_connections(29);
  `device_slave_connections(30);
  `device_slave_connections(31);
  `device_slave_connections(32);
  `device_slave_connections(33);
  `device_slave_connections(34);
  `device_slave_connections(35);
  `device_slave_connections(36);
  `device_slave_connections(37);
  `device_slave_connections(38);
  `device_slave_connections(39);
  `device_slave_connections(40);
  `device_slave_connections(41);
  `device_slave_connections(42);
  `device_slave_connections(43);
  `device_slave_connections(44);
  `device_slave_connections(45);
  `device_slave_connections(46);
  `device_slave_connections(47);
  `device_slave_connections(48);
  `device_slave_connections(49);
  `device_slave_connections(50);
  `device_slave_connections(51);
  `device_slave_connections(52);
  `device_slave_connections(53);
  `device_slave_connections(54);
  `device_slave_connections(55);
  `device_slave_connections(56);
  `device_slave_connections(57);
  `device_slave_connections(58);
  `device_slave_connections(59);
  `device_slave_connections(60);
  `device_slave_connections(61);
  `device_slave_connections(62);
  `device_slave_connections(63);
  `device_slave_connections(64);
  `device_slave_connections(65);
  `device_slave_connections(66);
  `device_slave_connections(67);
  `device_slave_connections(68);
  `device_slave_connections(69);
  `device_slave_connections(70);
  `device_slave_connections(71);
  `device_slave_connections(72);
  `device_slave_connections(73);
  `device_slave_connections(74);
  `device_slave_connections(75);
  `device_slave_connections(76);
  `device_slave_connections(77);
  `device_slave_connections(78);
  `device_slave_connections(79);
  `device_slave_connections(80);
  `device_slave_connections(81);
  `device_slave_connections(82);
  `device_slave_connections(83);
  `device_slave_connections(84);
  `device_slave_connections(85);
  `device_slave_connections(86);
  `device_slave_connections(87);
  `device_slave_connections(88);
  `device_slave_connections(89);
  `device_slave_connections(90);
  `device_slave_connections(91);
  `device_slave_connections(92);
  `device_slave_connections(93);
  `device_slave_connections(94);
  `device_slave_connections(95);
  `device_slave_connections(96);
  `device_slave_connections(97);
  `device_slave_connections(98);
  `device_slave_connections(99);
  `device_slave_connections(100);
  `device_slave_connections(101);
  `device_slave_connections(102);
  `device_slave_connections(103);
  `device_slave_connections(104);
  `device_slave_connections(105);
  `device_slave_connections(106);
  `device_slave_connections(107);
  `device_slave_connections(108);
  `device_slave_connections(109);
  `device_slave_connections(110);
  `device_slave_connections(111);
  `device_slave_connections(112);
  `device_slave_connections(113);
  `device_slave_connections(114);
  `device_slave_connections(115);
  `device_slave_connections(116);
  `device_slave_connections(117);
  `device_slave_connections(118);
  `device_slave_connections(119);
  `device_slave_connections(120);
  `device_slave_connections(121);
  `device_slave_connections(122);
  `device_slave_connections(123);
  `device_slave_connections(124);
  `device_slave_connections(125);
  `device_slave_connections(126);
  `device_slave_connections(127);
  `device_slave_connections(128);
  `device_slave_connections(129);
  `device_slave_connections(130);
  `device_slave_connections(131);
  `device_slave_connections(132);
  `device_slave_connections(133);
  `device_slave_connections(134);
  `device_slave_connections(135);
  `device_slave_connections(136);
  `device_slave_connections(137);
  `device_slave_connections(138);
  `device_slave_connections(139);
  `device_slave_connections(140);
  `device_slave_connections(141);
  `device_slave_connections(142);
  `device_slave_connections(143);
  `device_slave_connections(144);
  `device_slave_connections(145);
  `device_slave_connections(146);
  `device_slave_connections(147);
  `device_slave_connections(148);
  `device_slave_connections(149);
  `device_slave_connections(150);
  `device_slave_connections(151);
  `device_slave_connections(152);
  `device_slave_connections(153);
  `device_slave_connections(154);
  `device_slave_connections(155);
  `device_slave_connections(156);
  `device_slave_connections(157);
  `device_slave_connections(158);
  `device_slave_connections(159);
  `device_slave_connections(160);
  `device_slave_connections(161);
  `device_slave_connections(162);
  `device_slave_connections(163);
  `device_slave_connections(164);
  `device_slave_connections(165);
  `device_slave_connections(166);
  `device_slave_connections(167);
  `device_slave_connections(168);
  `device_slave_connections(169);
  `device_slave_connections(170);
  `device_slave_connections(171);
  `device_slave_connections(172);
  `device_slave_connections(173);
  `device_slave_connections(174);
  `device_slave_connections(175);
  `device_slave_connections(176);
  `device_slave_connections(177);
  `device_slave_connections(178);
  `device_slave_connections(179);
  `device_slave_connections(180);
  `device_slave_connections(181);
  `device_slave_connections(182);
  `device_slave_connections(183);
  `device_slave_connections(184);
  `device_slave_connections(185);
  `device_slave_connections(186);
  `device_slave_connections(187);
  `device_slave_connections(188);
  `device_slave_connections(189);
  `device_slave_connections(190);
  `device_slave_connections(191);
  `device_slave_connections(192);
  `device_slave_connections(193);
  `device_slave_connections(194);
  `device_slave_connections(195);
  `device_slave_connections(196);
  `device_slave_connections(197);
  `device_slave_connections(198);
  `device_slave_connections(199);
  `device_slave_connections(200);
  `device_slave_connections(201);
  `device_slave_connections(202);
  `device_slave_connections(203);
  `device_slave_connections(204);
  `device_slave_connections(205);
  `device_slave_connections(206);
  `device_slave_connections(207);
  `device_slave_connections(208);
  `device_slave_connections(209);
  `device_slave_connections(210);
  `device_slave_connections(211);
  `device_slave_connections(212);
  `device_slave_connections(213);
  `device_slave_connections(214);
  `device_slave_connections(215);
  `device_slave_connections(216);
  `device_slave_connections(217);
  `device_slave_connections(218);
  `device_slave_connections(219);
  `device_slave_connections(220);
  `device_slave_connections(221);
  `device_slave_connections(222);
  `device_slave_connections(223);
  `device_slave_connections(224);
  `device_slave_connections(225);
  `device_slave_connections(226);
  `device_slave_connections(227);
  `device_slave_connections(228);
  `device_slave_connections(229);
  `device_slave_connections(230);
  `device_slave_connections(231);
  `device_slave_connections(232);
  `device_slave_connections(233);
  `device_slave_connections(234);
  `device_slave_connections(235);
  `device_slave_connections(236);
  `device_slave_connections(237);
  `device_slave_connections(238);
  `device_slave_connections(239);
  `device_slave_connections(240);
  `device_slave_connections(241);
  `device_slave_connections(242);
  `device_slave_connections(243);
  `device_slave_connections(244);
  `device_slave_connections(245);
  `device_slave_connections(246);
  `device_slave_connections(247);
  `device_slave_connections(248);
  `device_slave_connections(249);
  `device_slave_connections(250);
  `device_slave_connections(251);
  `device_slave_connections(252);
  `device_slave_connections(253);
  `device_slave_connections(254);
  `device_slave_connections(255);
  `device_slave_connections(256);
  `device_slave_connections(257);
  `device_slave_connections(258);
  `device_slave_connections(259);
  `device_slave_connections(260);
  `device_slave_connections(261);
  `device_slave_connections(262);
  `device_slave_connections(263);
  `device_slave_connections(264);
  `device_slave_connections(265);
  `device_slave_connections(266);
  `device_slave_connections(267);
  `device_slave_connections(268);
  `device_slave_connections(269);
  `device_slave_connections(270);
  `device_slave_connections(271);
  `device_slave_connections(272);
  `device_slave_connections(273);
  `device_slave_connections(274);
  `device_slave_connections(275);
  `device_slave_connections(276);
  `device_slave_connections(277);
  `device_slave_connections(278);
  `device_slave_connections(279);
  `device_slave_connections(280);
  `device_slave_connections(281);
  `device_slave_connections(282);
  `device_slave_connections(283);
  `device_slave_connections(284);
  `device_slave_connections(285);
  `device_slave_connections(286);
  `device_slave_connections(287);
  `device_slave_connections(288);
  `device_slave_connections(289);
  `device_slave_connections(290);
  `device_slave_connections(291);
  `device_slave_connections(292);
  `device_slave_connections(293);
  `device_slave_connections(294);
  `device_slave_connections(295);
  `device_slave_connections(296);
  `device_slave_connections(297);
  `device_slave_connections(298);
  `device_slave_connections(299);
  `device_slave_connections(300);
  `device_slave_connections(301);
  `device_slave_connections(302);
  `device_slave_connections(303);
  `device_slave_connections(304);
  `device_slave_connections(305);
  `device_slave_connections(306);
  `device_slave_connections(307);
  `device_slave_connections(308);
  `device_slave_connections(309);
  `device_slave_connections(310);
  `device_slave_connections(311);
  `device_slave_connections(312);
  `device_slave_connections(313);
  `device_slave_connections(314);
  `device_slave_connections(315);
  `device_slave_connections(316);
  `device_slave_connections(317);
  `device_slave_connections(318);
  `device_slave_connections(319);
  `device_slave_connections(320);
  `device_slave_connections(321);
  `device_slave_connections(322);
  `device_slave_connections(323);
  `device_slave_connections(324);
  `device_slave_connections(325);
  `device_slave_connections(326);
  `device_slave_connections(327);
  `device_slave_connections(328);
  `device_slave_connections(329);
  `device_slave_connections(330);
  `device_slave_connections(331);
  `device_slave_connections(332);
  `device_slave_connections(333);
  `device_slave_connections(334);
  `device_slave_connections(335);
  `device_slave_connections(336);
  `device_slave_connections(337);
  `device_slave_connections(338);
  `device_slave_connections(339);
  `device_slave_connections(340);
  `device_slave_connections(341);
  `device_slave_connections(342);
  `device_slave_connections(343);
  `device_slave_connections(344);
  `device_slave_connections(345);
  `device_slave_connections(346);
  `device_slave_connections(347);
  `device_slave_connections(348);
  `device_slave_connections(349);
  `device_slave_connections(350);
  `device_slave_connections(351);
  `device_slave_connections(352);
  `device_slave_connections(353);
  `device_slave_connections(354);
  `device_slave_connections(355);
  `device_slave_connections(356);
  `device_slave_connections(357);
  `device_slave_connections(358);
  `device_slave_connections(359);
  `device_slave_connections(360);
  `device_slave_connections(361);
  `device_slave_connections(362);
  `device_slave_connections(363);
  `device_slave_connections(364);
  `device_slave_connections(365);
  `device_slave_connections(366);
  `device_slave_connections(367);
  `device_slave_connections(368);
  `device_slave_connections(369);
  `device_slave_connections(370);
  `device_slave_connections(371);
  `device_slave_connections(372);
  `device_slave_connections(373);
  `device_slave_connections(374);
  `device_slave_connections(375);
  `device_slave_connections(376);
  `device_slave_connections(377);
  `device_slave_connections(378);
  `device_slave_connections(379);
  `device_slave_connections(380);
  `device_slave_connections(381);
  `device_slave_connections(382);
  `device_slave_connections(383);
  `device_slave_connections(384);
  `device_slave_connections(385);
  `device_slave_connections(386);
  `device_slave_connections(387);
  `device_slave_connections(388);
  `device_slave_connections(389);
  `device_slave_connections(390);
  `device_slave_connections(391);
  `device_slave_connections(392);
  `device_slave_connections(393);
  `device_slave_connections(394);
  `device_slave_connections(395);
  `device_slave_connections(396);
  `device_slave_connections(397);
  `device_slave_connections(398);
  `device_slave_connections(399);
  `device_slave_connections(400);
  `device_slave_connections(401);
  `device_slave_connections(402);
  `device_slave_connections(403);
  `device_slave_connections(404);
  `device_slave_connections(405);
  `device_slave_connections(406);
  `device_slave_connections(407);
  `device_slave_connections(408);
  `device_slave_connections(409);
  `device_slave_connections(410);
  `device_slave_connections(411);
  `device_slave_connections(412);
  `device_slave_connections(413);
  `device_slave_connections(414);
  `device_slave_connections(415);
  `device_slave_connections(416);
  `device_slave_connections(417);
  `device_slave_connections(418);
  `device_slave_connections(419);
  `device_slave_connections(420);
  `device_slave_connections(421);
  `device_slave_connections(422);
  `device_slave_connections(423);
  `device_slave_connections(424);
  `device_slave_connections(425);
  `device_slave_connections(426);
  `device_slave_connections(427);
  `device_slave_connections(428);
  `device_slave_connections(429);
  `device_slave_connections(430);
  `device_slave_connections(431);
  `device_slave_connections(432);
  `device_slave_connections(433);
  `device_slave_connections(434);
  `device_slave_connections(435);
  `device_slave_connections(436);
  `device_slave_connections(437);
  `device_slave_connections(438);
  `device_slave_connections(439);
  `device_slave_connections(440);
  `device_slave_connections(441);
  `device_slave_connections(442);
  `device_slave_connections(443);
  `device_slave_connections(444);
  `device_slave_connections(445);
  `device_slave_connections(446);
  `device_slave_connections(447);
  `device_slave_connections(448);
  `device_slave_connections(449);
	`device_slave_connections_TB_CONFIG_4(0,450,0);
  `device_slave_connections_TB_CONFIG_4(0,451,1);
  `device_slave_connections_TB_CONFIG_4(0,452,2);
  `device_slave_connections_TB_CONFIG_4(0,453,3);
  `device_slave_connections_TB_CONFIG_4(0,454,4);
  `device_slave_connections_TB_CONFIG_4(0,455,5);
  `device_slave_connections_TB_CONFIG_4(0,456,6);
  `device_slave_connections_TB_CONFIG_4(0,457,7);
  `device_slave_connections_TB_CONFIG_4(0,458,8);
  `device_slave_connections_TB_CONFIG_4(0,459,9);
  `device_slave_connections_TB_CONFIG_4(0,460,10);
  `device_slave_connections_TB_CONFIG_4(0,461,11);
  `device_slave_connections_TB_CONFIG_4(0,462,12);
  `device_slave_connections_TB_CONFIG_4(0,463,13);
  `device_slave_connections_TB_CONFIG_4(0,464,14);
  `device_slave_connections_TB_CONFIG_4(0,465,15);
  `device_slave_connections_TB_CONFIG_4(0,466,16);
  `device_slave_connections_TB_CONFIG_4(0,467,17);
  `device_slave_connections_TB_CONFIG_4(0,468,18);
  `device_slave_connections_TB_CONFIG_4(0,469,19);
  `device_slave_connections_TB_CONFIG_4(0,470,20);
  `device_slave_connections_TB_CONFIG_4(0,471,21);
  `device_slave_connections_TB_CONFIG_4(0,472,22);
  `device_slave_connections_TB_CONFIG_4(0,473,23);
  `device_slave_connections_TB_CONFIG_4(0,474,24);
  `device_slave_connections_TB_CONFIG_4(0,475,25);
  `device_slave_connections_TB_CONFIG_4(0,476,26);
  `device_slave_connections_TB_CONFIG_4(0,477,27);
  `device_slave_connections_TB_CONFIG_4(0,478,28);
  `device_slave_connections_TB_CONFIG_4(0,479,29);
  `device_slave_connections_TB_CONFIG_4(0,480,30);
  `device_slave_connections_TB_CONFIG_4(0,481,31);
  `device_slave_connections_TB_CONFIG_4(0,482,32);
  `device_slave_connections_TB_CONFIG_4(0,483,33);
  `device_slave_connections_TB_CONFIG_4(0,484,34);
  `device_slave_connections_TB_CONFIG_4(0,485,35);
  `device_slave_connections_TB_CONFIG_4(0,486,36);
  `device_slave_connections_TB_CONFIG_4(0,487,37);
  `device_slave_connections_TB_CONFIG_4(0,488,38);
  `device_slave_connections_TB_CONFIG_4(0,489,39);
  `device_slave_connections_TB_CONFIG_4(0,490,40);
  `device_slave_connections_TB_CONFIG_4(0,491,41);
  `device_slave_connections_TB_CONFIG_4(0,492,42);
  `device_slave_connections_TB_CONFIG_4(0,493,43);
  `device_slave_connections_TB_CONFIG_4(0,494,44);
  `device_slave_connections_TB_CONFIG_4(0,495,45);
  `device_slave_connections_TB_CONFIG_4(0,496,46);
  `device_slave_connections_TB_CONFIG_4(0,497,47);
  `device_slave_connections_TB_CONFIG_4(0,498,48);
  `device_slave_connections_TB_CONFIG_4(0,499,49);
  `device_slave_connections_TB_CONFIG_4(0,500,50);
  `device_slave_connections_TB_CONFIG_4(0,501,51);
  `device_slave_connections_TB_CONFIG_4(0,502,52);
  `device_slave_connections_TB_CONFIG_4(0,503,53);
  `device_slave_connections_TB_CONFIG_4(0,504,54);
  `device_slave_connections_TB_CONFIG_4(0,505,55);
  `device_slave_connections_TB_CONFIG_4(0,506,56);
  `device_slave_connections_TB_CONFIG_4(0,507,57);
  `device_slave_connections_TB_CONFIG_4(0,508,58);
  `device_slave_connections_TB_CONFIG_4(0,509,59);
  `device_slave_connections_TB_CONFIG_4(0,510,60);
  `device_slave_connections_TB_CONFIG_4(0,511,61);
  `device_slave_connections_TB_CONFIG_4(0,512,62);
  `device_slave_connections_TB_CONFIG_4(0,513,63);
  `device_slave_connections_TB_CONFIG_4(0,514,64);
  `device_slave_connections_TB_CONFIG_4(0,515,65);
  `device_slave_connections_TB_CONFIG_4(0,516,66);
  `device_slave_connections_TB_CONFIG_4(0,517,67);
  `device_slave_connections_TB_CONFIG_4(0,518,68);
  `device_slave_connections_TB_CONFIG_4(0,519,69);
  `device_slave_connections_TB_CONFIG_4(0,520,70);
  `device_slave_connections_TB_CONFIG_4(0,521,71);
  `device_slave_connections_TB_CONFIG_4(0,522,72);
  `device_slave_connections_TB_CONFIG_4(0,523,73);
  `device_slave_connections_TB_CONFIG_4(0,524,74);
  `device_slave_connections_TB_CONFIG_4(0,525,75);
  `device_slave_connections_TB_CONFIG_4(0,526,76);
  `device_slave_connections_TB_CONFIG_4(0,527,77);
  `device_slave_connections_TB_CONFIG_4(0,528,78);
  `device_slave_connections_TB_CONFIG_4(0,529,79);
  `device_slave_connections_TB_CONFIG_4(0,530,80);
  `device_slave_connections_TB_CONFIG_4(0,531,81);
  `device_slave_connections_TB_CONFIG_4(0,532,82);
  `device_slave_connections_TB_CONFIG_4(0,533,83);
  `device_slave_connections_TB_CONFIG_4(0,534,84);
  `device_slave_connections_TB_CONFIG_4(0,535,85);
  `device_slave_connections_TB_CONFIG_4(0,536,86);
  `device_slave_connections_TB_CONFIG_4(0,537,87);
  `device_slave_connections_TB_CONFIG_4(0,538,88);
  `device_slave_connections_TB_CONFIG_4(0,539,89);
  `device_slave_connections_TB_CONFIG_4(0,540,90);
  `device_slave_connections_TB_CONFIG_4(0,541,91);
  `device_slave_connections_TB_CONFIG_4(0,542,92);
  `device_slave_connections_TB_CONFIG_4(0,543,93);
  `device_slave_connections_TB_CONFIG_4(0,544,94);
  `device_slave_connections_TB_CONFIG_4(0,545,95);
  `device_slave_connections_TB_CONFIG_4(0,546,96);
  `device_slave_connections_TB_CONFIG_4(0,547,97);
  `device_slave_connections_TB_CONFIG_4(0,548,98);
  `device_slave_connections_TB_CONFIG_4(0,549,99);
  `device_slave_connections_TB_CONFIG_4(0,550,100);
  `device_slave_connections_TB_CONFIG_4(0,551,101);
  `device_slave_connections_TB_CONFIG_4(0,552,102);
  `device_slave_connections_TB_CONFIG_4(0,553,103);
  `device_slave_connections_TB_CONFIG_4(0,554,104);
  `device_slave_connections_TB_CONFIG_4(0,555,105);
  `device_slave_connections_TB_CONFIG_4(0,556,106);
  `device_slave_connections_TB_CONFIG_4(0,557,107);
  `device_slave_connections_TB_CONFIG_4(0,558,108);
  `device_slave_connections_TB_CONFIG_4(0,559,109);
  `device_slave_connections_TB_CONFIG_4(0,560,110);
  `device_slave_connections_TB_CONFIG_4(0,561,111);
  `device_slave_connections_TB_CONFIG_4(0,562,112);
  `device_slave_connections_TB_CONFIG_4(0,563,113);
  `device_slave_connections_TB_CONFIG_4(0,564,114);
  `device_slave_connections_TB_CONFIG_4(0,565,115);
  `device_slave_connections_TB_CONFIG_4(0,566,116);
  `device_slave_connections_TB_CONFIG_4(0,567,117);
  `device_slave_connections_TB_CONFIG_4(0,568,118);
  `device_slave_connections_TB_CONFIG_4(0,569,119);
  `device_slave_connections_TB_CONFIG_4(0,570,120);
  `device_slave_connections_TB_CONFIG_4(0,571,121);
  `device_slave_connections_TB_CONFIG_4(0,572,122);
  `device_slave_connections_TB_CONFIG_4(0,573,123);
  `device_slave_connections_TB_CONFIG_4(0,574,124);
  `device_slave_connections_TB_CONFIG_4(0,575,125);
  `device_slave_connections_TB_CONFIG_4(0,576,126);
  `device_slave_connections_TB_CONFIG_4(0,577,127);
  `device_slave_connections_TB_CONFIG_4(0,578,128);
  `device_slave_connections_TB_CONFIG_4(0,579,129);
  `device_slave_connections_TB_CONFIG_4(0,580,130);
  `device_slave_connections_TB_CONFIG_4(0,581,131);
  `device_slave_connections_TB_CONFIG_4(0,582,132);
  `device_slave_connections_TB_CONFIG_4(0,583,133);
  `device_slave_connections_TB_CONFIG_4(0,584,134);
  `device_slave_connections_TB_CONFIG_4(0,585,135);
  `device_slave_connections_TB_CONFIG_4(0,586,136);
  `device_slave_connections_TB_CONFIG_4(0,587,137);
  `device_slave_connections_TB_CONFIG_4(0,588,138);
  `device_slave_connections_TB_CONFIG_4(0,589,139);
  `device_slave_connections_TB_CONFIG_4(0,590,140);
  `device_slave_connections_TB_CONFIG_4(0,591,141);
  `device_slave_connections_TB_CONFIG_4(0,592,142);
  `device_slave_connections_TB_CONFIG_4(0,593,143);
  `device_slave_connections_TB_CONFIG_4(0,594,144);
  `device_slave_connections_TB_CONFIG_4(0,595,145);
  `device_slave_connections_TB_CONFIG_4(0,596,146);
  `device_slave_connections_TB_CONFIG_4(0,597,147);
  `device_slave_connections_TB_CONFIG_4(0,598,148);
  `device_slave_connections_TB_CONFIG_4(0,599,149);
  `device_slave_connections_TB_CONFIG_4(0,600,150);
  `device_slave_connections_TB_CONFIG_4(0,601,151);
  `device_slave_connections_TB_CONFIG_4(0,602,152);
  `device_slave_connections_TB_CONFIG_4(0,603,153);
  `device_slave_connections_TB_CONFIG_4(0,604,154);
  `device_slave_connections_TB_CONFIG_4(0,605,155);
  `device_slave_connections_TB_CONFIG_4(0,606,156);
  `device_slave_connections_TB_CONFIG_4(0,607,157);
  `device_slave_connections_TB_CONFIG_4(0,608,158);
  `device_slave_connections_TB_CONFIG_4(0,609,159);
  `device_slave_connections_TB_CONFIG_4(0,610,160);
  `device_slave_connections_TB_CONFIG_4(0,611,161);
  `device_slave_connections_TB_CONFIG_4(0,612,162);
  `device_slave_connections_TB_CONFIG_4(0,613,163);
  `device_slave_connections_TB_CONFIG_4(0,614,164);
  `device_slave_connections_TB_CONFIG_4(0,615,165);
  `device_slave_connections_TB_CONFIG_4(0,616,166);
  `device_slave_connections_TB_CONFIG_4(0,617,167);
  `device_slave_connections_TB_CONFIG_4(0,618,168);
  `device_slave_connections_TB_CONFIG_4(0,619,169);
  `device_slave_connections_TB_CONFIG_4(0,620,170);
  `device_slave_connections_TB_CONFIG_4(0,621,171);
  `device_slave_connections_TB_CONFIG_4(0,622,172);
  `device_slave_connections_TB_CONFIG_4(0,623,173);
  `device_slave_connections_TB_CONFIG_4(0,624,174);
  `device_slave_connections_TB_CONFIG_4(0,625,175);
  `device_slave_connections_TB_CONFIG_4(0,626,176);
  `device_slave_connections_TB_CONFIG_4(0,627,177);
  `device_slave_connections_TB_CONFIG_4(0,628,178);
  `device_slave_connections_TB_CONFIG_4(0,629,179);
  `device_slave_connections_TB_CONFIG_4(0,630,180);
  `device_slave_connections_TB_CONFIG_4(0,631,181);
  `device_slave_connections_TB_CONFIG_4(0,632,182);
  `device_slave_connections_TB_CONFIG_4(0,633,183);
  `device_slave_connections_TB_CONFIG_4(0,634,184);
  `device_slave_connections_TB_CONFIG_4(0,635,185);
  `device_slave_connections_TB_CONFIG_4(0,636,186);
  `device_slave_connections_TB_CONFIG_4(0,637,187);
  `device_slave_connections_TB_CONFIG_4(0,638,188);
  `device_slave_connections_TB_CONFIG_4(0,639,189);
  `device_slave_connections_TB_CONFIG_4(0,640,190);
  `device_slave_connections_TB_CONFIG_4(0,641,191);
  `device_slave_connections_TB_CONFIG_4(0,642,192);
  `device_slave_connections_TB_CONFIG_4(0,643,193);
  `device_slave_connections_TB_CONFIG_4(0,644,194);
  `device_slave_connections_TB_CONFIG_4(0,645,195);
  `device_slave_connections_TB_CONFIG_4(0,646,196);
  `device_slave_connections_TB_CONFIG_4(0,647,197);
  `device_slave_connections_TB_CONFIG_4(0,648,198);
  `device_slave_connections_TB_CONFIG_4(0,649,199);
  `device_slave_connections_TB_CONFIG_4(0,650,200);
  `device_slave_connections_TB_CONFIG_4(0,651,201);
  `device_slave_connections_TB_CONFIG_4(0,652,202);
  `device_slave_connections_TB_CONFIG_4(0,653,203);
  `device_slave_connections_TB_CONFIG_4(0,654,204);
  `device_slave_connections_TB_CONFIG_4(0,655,205);
  `device_slave_connections_TB_CONFIG_4(0,656,206);
  `device_slave_connections_TB_CONFIG_4(0,657,207);
  `device_slave_connections_TB_CONFIG_4(0,658,208);
  `device_slave_connections_TB_CONFIG_4(0,659,209);
  `device_slave_connections_TB_CONFIG_4(0,660,210);
  `device_slave_connections_TB_CONFIG_4(0,661,211);
  `device_slave_connections_TB_CONFIG_4(0,662,212);
  `device_slave_connections_TB_CONFIG_4(0,663,213);
  `device_slave_connections_TB_CONFIG_4(0,664,214);
  `device_slave_connections_TB_CONFIG_4(0,665,215);
  `device_slave_connections_TB_CONFIG_4(0,666,216);
  `device_slave_connections_TB_CONFIG_4(0,667,217);
  `device_slave_connections_TB_CONFIG_4(0,668,218);
  `device_slave_connections_TB_CONFIG_4(0,669,219);
  `device_slave_connections_TB_CONFIG_4(0,670,220);
  `device_slave_connections_TB_CONFIG_4(0,671,221);
  `device_slave_connections_TB_CONFIG_4(0,672,222);
  `device_slave_connections_TB_CONFIG_4(0,673,223);
  `device_slave_connections_TB_CONFIG_4(0,674,224);
  `device_slave_connections_TB_CONFIG_4(0,675,225);
  `device_slave_connections_TB_CONFIG_4(0,676,226);
  `device_slave_connections_TB_CONFIG_4(0,677,227);
  `device_slave_connections_TB_CONFIG_4(0,678,228);
  `device_slave_connections_TB_CONFIG_4(0,679,229);
  `device_slave_connections_TB_CONFIG_4(0,680,230);
  `device_slave_connections_TB_CONFIG_4(0,681,231);
  `device_slave_connections_TB_CONFIG_4(0,682,232);
  `device_slave_connections_TB_CONFIG_4(0,683,233);
  `device_slave_connections_TB_CONFIG_4(0,684,234);
  `device_slave_connections_TB_CONFIG_4(0,685,235);
  `device_slave_connections_TB_CONFIG_4(0,686,236);
  `device_slave_connections_TB_CONFIG_4(0,687,237);
  `device_slave_connections_TB_CONFIG_4(0,688,238);
  `device_slave_connections_TB_CONFIG_4(0,689,239);
  `device_slave_connections_TB_CONFIG_4(0,690,240);
  `device_slave_connections_TB_CONFIG_4(0,691,241);
  `device_slave_connections_TB_CONFIG_4(0,692,242);
  `device_slave_connections_TB_CONFIG_4(0,693,243);
  `device_slave_connections_TB_CONFIG_4(0,694,244);
  `device_slave_connections_TB_CONFIG_4(0,695,245);
  `device_slave_connections_TB_CONFIG_4(0,696,246);
  `device_slave_connections_TB_CONFIG_4(0,697,247);
  `device_slave_connections_TB_CONFIG_4(0,698,248);
  `device_slave_connections_TB_CONFIG_4(0,699,249);
  `device_slave_connections_TB_CONFIG_4(0,700,250);
  `device_slave_connections_TB_CONFIG_4(0,701,251);
  `device_slave_connections_TB_CONFIG_4(0,702,252);
  `device_slave_connections_TB_CONFIG_4(0,703,253);
  `device_slave_connections_TB_CONFIG_4(0,704,254);
  `device_slave_connections_TB_CONFIG_4(0,705,255);
  `device_slave_connections_TB_CONFIG_4(0,706,256);
  `device_slave_connections_TB_CONFIG_4(0,707,257);
  `device_slave_connections_TB_CONFIG_4(0,708,258);
  `device_slave_connections_TB_CONFIG_4(0,709,259);
  `device_slave_connections_TB_CONFIG_4(0,710,260);
  `device_slave_connections_TB_CONFIG_4(0,711,261);
  `device_slave_connections_TB_CONFIG_4(0,712,262);
  `device_slave_connections_TB_CONFIG_4(0,713,263);
  `device_slave_connections_TB_CONFIG_4(0,714,264);
  `device_slave_connections_TB_CONFIG_4(0,715,265);
  `device_slave_connections_TB_CONFIG_4(0,716,266);
  `device_slave_connections_TB_CONFIG_4(0,717,267);
  `device_slave_connections_TB_CONFIG_4(0,718,268);
  `device_slave_connections_TB_CONFIG_4(0,719,269);
  `device_slave_connections_TB_CONFIG_4(0,720,270);
  `device_slave_connections_TB_CONFIG_4(0,721,271);
  `device_slave_connections_TB_CONFIG_4(0,722,272);
  `device_slave_connections_TB_CONFIG_4(0,723,273);
  `device_slave_connections_TB_CONFIG_4(0,724,274);
  `device_slave_connections_TB_CONFIG_4(0,725,275);
  `device_slave_connections_TB_CONFIG_4(0,726,276);
  `device_slave_connections_TB_CONFIG_4(0,727,277);
  `device_slave_connections_TB_CONFIG_4(0,728,278);
  `device_slave_connections_TB_CONFIG_4(0,729,279);
  `device_slave_connections_TB_CONFIG_4(0,730,280);
  `device_slave_connections_TB_CONFIG_4(0,731,281);
  `device_slave_connections_TB_CONFIG_4(0,732,282);
  `device_slave_connections_TB_CONFIG_4(0,733,283);
  `device_slave_connections_TB_CONFIG_4(0,734,284);
  `device_slave_connections_TB_CONFIG_4(0,735,285);
  `device_slave_connections_TB_CONFIG_4(0,736,286);
  `device_slave_connections_TB_CONFIG_4(0,737,287);
  `device_slave_connections_TB_CONFIG_4(0,738,288);
  `device_slave_connections_TB_CONFIG_4(0,739,289);
  `device_slave_connections_TB_CONFIG_4(0,740,290);
  `device_slave_connections_TB_CONFIG_4(0,741,291);
  `device_slave_connections_TB_CONFIG_4(0,742,292);
  `device_slave_connections_TB_CONFIG_4(0,743,293);
  `device_slave_connections_TB_CONFIG_4(0,744,294);
  `device_slave_connections_TB_CONFIG_4(0,745,295);
  `device_slave_connections_TB_CONFIG_4(0,746,296);
  `device_slave_connections_TB_CONFIG_4(0,747,297);
  `device_slave_connections_TB_CONFIG_4(0,748,298);
  `device_slave_connections_TB_CONFIG_4(0,749,299);
  `device_slave_connections_TB_CONFIG_4(0,750,300);
  `device_slave_connections_TB_CONFIG_4(0,751,301);
  `device_slave_connections_TB_CONFIG_4(0,752,302);
  `device_slave_connections_TB_CONFIG_4(0,753,303);
  `device_slave_connections_TB_CONFIG_4(0,754,304);
  `device_slave_connections_TB_CONFIG_4(0,755,305);
  `device_slave_connections_TB_CONFIG_4(0,756,306);
  `device_slave_connections_TB_CONFIG_4(0,757,307);
  `device_slave_connections_TB_CONFIG_4(0,758,308);
  `device_slave_connections_TB_CONFIG_4(0,759,309);
  `device_slave_connections_TB_CONFIG_4(0,760,310);
  `device_slave_connections_TB_CONFIG_4(0,761,311);
  `device_slave_connections_TB_CONFIG_4(0,762,312);
  `device_slave_connections_TB_CONFIG_4(0,763,313);
  `device_slave_connections_TB_CONFIG_4(0,764,314);
  `device_slave_connections_TB_CONFIG_4(0,765,315);
  `device_slave_connections_TB_CONFIG_4(0,766,316);
  `device_slave_connections_TB_CONFIG_4(0,767,317);
  `device_slave_connections_TB_CONFIG_4(0,768,318);
  `device_slave_connections_TB_CONFIG_4(0,769,319);
  `device_slave_connections_TB_CONFIG_4(0,770,320);
  `device_slave_connections_TB_CONFIG_4(0,771,321);
  `device_slave_connections_TB_CONFIG_4(0,772,322);
  `device_slave_connections_TB_CONFIG_4(0,773,323);
  `device_slave_connections_TB_CONFIG_4(0,774,324);
  `device_slave_connections_TB_CONFIG_4(0,775,325);
  `device_slave_connections_TB_CONFIG_4(0,776,326);
  `device_slave_connections_TB_CONFIG_4(0,777,327);
  `device_slave_connections_TB_CONFIG_4(0,778,328);
  `device_slave_connections_TB_CONFIG_4(0,779,329);
  `device_slave_connections_TB_CONFIG_4(0,780,330);
  `device_slave_connections_TB_CONFIG_4(0,781,331);
  `device_slave_connections_TB_CONFIG_4(0,782,332);
  `device_slave_connections_TB_CONFIG_4(0,783,333);
  `device_slave_connections_TB_CONFIG_4(0,784,334);
  `device_slave_connections_TB_CONFIG_4(0,785,335);
  `device_slave_connections_TB_CONFIG_4(0,786,336);
  `device_slave_connections_TB_CONFIG_4(0,787,337);
  `device_slave_connections_TB_CONFIG_4(0,788,338);
  `device_slave_connections_TB_CONFIG_4(0,789,339);
  `device_slave_connections_TB_CONFIG_4(0,790,340);
  `device_slave_connections_TB_CONFIG_4(0,791,341);
  `device_slave_connections_TB_CONFIG_4(0,792,342);
  `device_slave_connections_TB_CONFIG_4(0,793,343);
  `device_slave_connections_TB_CONFIG_4(0,794,344);
  `device_slave_connections_TB_CONFIG_4(0,795,345);
  `device_slave_connections_TB_CONFIG_4(0,796,346);
  `device_slave_connections_TB_CONFIG_4(0,797,347);
  `device_slave_connections_TB_CONFIG_4(0,798,348);
  `device_slave_connections_TB_CONFIG_4(0,799,349);
  `device_slave_connections_TB_CONFIG_4(0,800,350);
  `device_slave_connections_TB_CONFIG_4(0,801,351);
  `device_slave_connections_TB_CONFIG_4(0,802,352);
  `device_slave_connections_TB_CONFIG_4(0,803,353);
  `device_slave_connections_TB_CONFIG_4(0,804,354);
  `device_slave_connections_TB_CONFIG_4(0,805,355);
  `device_slave_connections_TB_CONFIG_4(0,806,356);
  `device_slave_connections_TB_CONFIG_4(0,807,357);
  `device_slave_connections_TB_CONFIG_4(0,808,358);
  `device_slave_connections_TB_CONFIG_4(0,809,359);
  `device_slave_connections_TB_CONFIG_4(0,810,360);
  `device_slave_connections_TB_CONFIG_4(0,811,361);
  `device_slave_connections_TB_CONFIG_4(0,812,362);
  `device_slave_connections_TB_CONFIG_4(0,813,363);
  `device_slave_connections_TB_CONFIG_4(0,814,364);
  `device_slave_connections_TB_CONFIG_4(0,815,365);
  `device_slave_connections_TB_CONFIG_4(0,816,366);
  `device_slave_connections_TB_CONFIG_4(0,817,367);
  `device_slave_connections_TB_CONFIG_4(0,818,368);
  `device_slave_connections_TB_CONFIG_4(0,819,369);
  `device_slave_connections_TB_CONFIG_4(0,820,370);
  `device_slave_connections_TB_CONFIG_4(0,821,371);
  `device_slave_connections_TB_CONFIG_4(0,822,372);
  `device_slave_connections_TB_CONFIG_4(0,823,373);
  `device_slave_connections_TB_CONFIG_4(0,824,374);
  `device_slave_connections_TB_CONFIG_4(0,825,375);
  `device_slave_connections_TB_CONFIG_4(0,826,376);
  `device_slave_connections_TB_CONFIG_4(0,827,377);
  `device_slave_connections_TB_CONFIG_4(0,828,378);
  `device_slave_connections_TB_CONFIG_4(0,829,379);
  `device_slave_connections_TB_CONFIG_4(0,830,380);
  `device_slave_connections_TB_CONFIG_4(0,831,381);
  `device_slave_connections_TB_CONFIG_4(0,832,382);
  `device_slave_connections_TB_CONFIG_4(0,833,383);
  `device_slave_connections_TB_CONFIG_4(0,834,384);
  `device_slave_connections_TB_CONFIG_4(0,835,385);
  `device_slave_connections_TB_CONFIG_4(0,836,386);
  `device_slave_connections_TB_CONFIG_4(0,837,387);
  `device_slave_connections_TB_CONFIG_4(0,838,388);
  `device_slave_connections_TB_CONFIG_4(0,839,389);
  `device_slave_connections_TB_CONFIG_4(0,840,390);
  `device_slave_connections_TB_CONFIG_4(0,841,391);
  `device_slave_connections_TB_CONFIG_4(0,842,392);
  `device_slave_connections_TB_CONFIG_4(0,843,393);
  `device_slave_connections_TB_CONFIG_4(0,844,394);
  `device_slave_connections_TB_CONFIG_4(0,845,395);
  `device_slave_connections_TB_CONFIG_4(0,846,396);
  `device_slave_connections_TB_CONFIG_4(0,847,397);
  `device_slave_connections_TB_CONFIG_4(0,848,398);
  `device_slave_connections_TB_CONFIG_4(0,849,399);
  `device_slave_connections_TB_CONFIG_4(0,850,400);
  `device_slave_connections_TB_CONFIG_4(0,851,401);
  `device_slave_connections_TB_CONFIG_4(0,852,402);
  `device_slave_connections_TB_CONFIG_4(0,853,403);
  `device_slave_connections_TB_CONFIG_4(0,854,404);
  `device_slave_connections_TB_CONFIG_4(0,855,405);
  `device_slave_connections_TB_CONFIG_4(0,856,406);
  `device_slave_connections_TB_CONFIG_4(0,857,407);
  `device_slave_connections_TB_CONFIG_4(0,858,408);
  `device_slave_connections_TB_CONFIG_4(0,859,409);
  `device_slave_connections_TB_CONFIG_4(0,860,410);
  `device_slave_connections_TB_CONFIG_4(0,861,411);
  `device_slave_connections_TB_CONFIG_4(0,862,412);
  `device_slave_connections_TB_CONFIG_4(0,863,413);
  `device_slave_connections_TB_CONFIG_4(0,864,414);
  `device_slave_connections_TB_CONFIG_4(0,865,415);
  `device_slave_connections_TB_CONFIG_4(0,866,416);
  `device_slave_connections_TB_CONFIG_4(0,867,417);
  `device_slave_connections_TB_CONFIG_4(0,868,418);
  `device_slave_connections_TB_CONFIG_4(0,869,419);
  `device_slave_connections_TB_CONFIG_4(0,870,420);
  `device_slave_connections_TB_CONFIG_4(0,871,421);
  `device_slave_connections_TB_CONFIG_4(0,872,422);
  `device_slave_connections_TB_CONFIG_4(0,873,423);
  `device_slave_connections_TB_CONFIG_4(0,874,424);
  `device_slave_connections_TB_CONFIG_4(0,875,425);
  `device_slave_connections_TB_CONFIG_4(0,876,426);
  `device_slave_connections_TB_CONFIG_4(0,877,427);
  `device_slave_connections_TB_CONFIG_4(0,878,428);
  `device_slave_connections_TB_CONFIG_4(0,879,429);
  `device_slave_connections_TB_CONFIG_4(0,880,430);
  `device_slave_connections_TB_CONFIG_4(0,881,431);
  `device_slave_connections_TB_CONFIG_4(0,882,432);
  `device_slave_connections_TB_CONFIG_4(0,883,433);
  `device_slave_connections_TB_CONFIG_4(0,884,434);
  `device_slave_connections_TB_CONFIG_4(0,885,435);
  `device_slave_connections_TB_CONFIG_4(0,886,436);
  `device_slave_connections_TB_CONFIG_4(0,887,437);
  `device_slave_connections_TB_CONFIG_4(0,888,438);
  `device_slave_connections_TB_CONFIG_4(0,889,439);
  `device_slave_connections_TB_CONFIG_4(0,890,440);
  `device_slave_connections_TB_CONFIG_4(0,891,441);
  `device_slave_connections_TB_CONFIG_4(0,892,442);
  `device_slave_connections_TB_CONFIG_4(0,893,443);
  `device_slave_connections_TB_CONFIG_4(0,894,444);
  `device_slave_connections_TB_CONFIG_4(0,895,445);
  `device_slave_connections_TB_CONFIG_4(0,896,446);
  `device_slave_connections_TB_CONFIG_4(0,897,447);
  `device_slave_connections_TB_CONFIG_4(0,898,448);
  `device_slave_connections_TB_CONFIG_4(0,899,449);
  `device_slave_connections_TB_CONFIG_4(1,900,0);
  `device_slave_connections_TB_CONFIG_4(1,901,1);
  `device_slave_connections_TB_CONFIG_4(1,902,2);
  `device_slave_connections_TB_CONFIG_4(1,903,3);
  `device_slave_connections_TB_CONFIG_4(1,904,4);
  `device_slave_connections_TB_CONFIG_4(1,905,5);
  `device_slave_connections_TB_CONFIG_4(1,906,6);
  `device_slave_connections_TB_CONFIG_4(1,907,7);
  `device_slave_connections_TB_CONFIG_4(1,908,8);
  `device_slave_connections_TB_CONFIG_4(1,909,9);
  `device_slave_connections_TB_CONFIG_4(1,910,10);
  `device_slave_connections_TB_CONFIG_4(1,911,11);
  `device_slave_connections_TB_CONFIG_4(1,912,12);
  `device_slave_connections_TB_CONFIG_4(1,913,13);
  `device_slave_connections_TB_CONFIG_4(1,914,14);
  `device_slave_connections_TB_CONFIG_4(1,915,15);
  `device_slave_connections_TB_CONFIG_4(1,916,16);
  `device_slave_connections_TB_CONFIG_4(1,917,17);
  `device_slave_connections_TB_CONFIG_4(1,918,18);
  `device_slave_connections_TB_CONFIG_4(1,919,19);
  `device_slave_connections_TB_CONFIG_4(1,920,20);
  `device_slave_connections_TB_CONFIG_4(1,921,21);
  `device_slave_connections_TB_CONFIG_4(1,922,22);
  `device_slave_connections_TB_CONFIG_4(1,923,23);
  `device_slave_connections_TB_CONFIG_4(1,924,24);
  `device_slave_connections_TB_CONFIG_4(1,925,25);
  `device_slave_connections_TB_CONFIG_4(1,926,26);
  `device_slave_connections_TB_CONFIG_4(1,927,27);
  `device_slave_connections_TB_CONFIG_4(1,928,28);
  `device_slave_connections_TB_CONFIG_4(1,929,29);
  `device_slave_connections_TB_CONFIG_4(1,930,30);
  `device_slave_connections_TB_CONFIG_4(1,931,31);
  `device_slave_connections_TB_CONFIG_4(1,932,32);
  `device_slave_connections_TB_CONFIG_4(1,933,33);
  `device_slave_connections_TB_CONFIG_4(1,934,34);
  `device_slave_connections_TB_CONFIG_4(1,935,35);
  `device_slave_connections_TB_CONFIG_4(1,936,36);
  `device_slave_connections_TB_CONFIG_4(1,937,37);
  `device_slave_connections_TB_CONFIG_4(1,938,38);
  `device_slave_connections_TB_CONFIG_4(1,939,39);
  `device_slave_connections_TB_CONFIG_4(1,940,40);
  `device_slave_connections_TB_CONFIG_4(1,941,41);
  `device_slave_connections_TB_CONFIG_4(1,942,42);
  `device_slave_connections_TB_CONFIG_4(1,943,43);
  `device_slave_connections_TB_CONFIG_4(1,944,44);
  `device_slave_connections_TB_CONFIG_4(1,945,45);
  `device_slave_connections_TB_CONFIG_4(1,946,46);
  `device_slave_connections_TB_CONFIG_4(1,947,47);
  `device_slave_connections_TB_CONFIG_4(1,948,48);
  `device_slave_connections_TB_CONFIG_4(1,949,49);
  `device_slave_connections_TB_CONFIG_4(1,950,50);
  `device_slave_connections_TB_CONFIG_4(1,951,51);
  `device_slave_connections_TB_CONFIG_4(1,952,52);
  `device_slave_connections_TB_CONFIG_4(1,953,53);
  `device_slave_connections_TB_CONFIG_4(1,954,54);
  `device_slave_connections_TB_CONFIG_4(1,955,55);
  `device_slave_connections_TB_CONFIG_4(1,956,56);
  `device_slave_connections_TB_CONFIG_4(1,957,57);
  `device_slave_connections_TB_CONFIG_4(1,958,58);
  `device_slave_connections_TB_CONFIG_4(1,959,59);
  `device_slave_connections_TB_CONFIG_4(1,960,60);
  `device_slave_connections_TB_CONFIG_4(1,961,61);
  `device_slave_connections_TB_CONFIG_4(1,962,62);
  `device_slave_connections_TB_CONFIG_4(1,963,63);
  `device_slave_connections_TB_CONFIG_4(1,964,64);
  `device_slave_connections_TB_CONFIG_4(1,965,65);
  `device_slave_connections_TB_CONFIG_4(1,966,66);
  `device_slave_connections_TB_CONFIG_4(1,967,67);
  `device_slave_connections_TB_CONFIG_4(1,968,68);
  `device_slave_connections_TB_CONFIG_4(1,969,69);
  `device_slave_connections_TB_CONFIG_4(1,970,70);
  `device_slave_connections_TB_CONFIG_4(1,971,71);
  `device_slave_connections_TB_CONFIG_4(1,972,72);
  `device_slave_connections_TB_CONFIG_4(1,973,73);
  `device_slave_connections_TB_CONFIG_4(1,974,74);
  `device_slave_connections_TB_CONFIG_4(1,975,75);
  `device_slave_connections_TB_CONFIG_4(1,976,76);
  `device_slave_connections_TB_CONFIG_4(1,977,77);
  `device_slave_connections_TB_CONFIG_4(1,978,78);
  `device_slave_connections_TB_CONFIG_4(1,979,79);
  `device_slave_connections_TB_CONFIG_4(1,980,80);
  `device_slave_connections_TB_CONFIG_4(1,981,81);
  `device_slave_connections_TB_CONFIG_4(1,982,82);
  `device_slave_connections_TB_CONFIG_4(1,983,83);
  `device_slave_connections_TB_CONFIG_4(1,984,84);
  `device_slave_connections_TB_CONFIG_4(1,985,85);
  `device_slave_connections_TB_CONFIG_4(1,986,86);
  `device_slave_connections_TB_CONFIG_4(1,987,87);
  `device_slave_connections_TB_CONFIG_4(1,988,88);
  `device_slave_connections_TB_CONFIG_4(1,989,89);
  `device_slave_connections_TB_CONFIG_4(1,990,90);
  `device_slave_connections_TB_CONFIG_4(1,991,91);
  `device_slave_connections_TB_CONFIG_4(1,992,92);
  `device_slave_connections_TB_CONFIG_4(1,993,93);
  `device_slave_connections_TB_CONFIG_4(1,994,94);
  `device_slave_connections_TB_CONFIG_4(1,995,95);
  `device_slave_connections_TB_CONFIG_4(1,996,96);
  `device_slave_connections_TB_CONFIG_4(1,997,97);
  `device_slave_connections_TB_CONFIG_4(1,998,98);
  `device_slave_connections_TB_CONFIG_4(1,999,99);
  `device_slave_connections_TB_CONFIG_4(1,1000,100);
  `device_slave_connections_TB_CONFIG_4(1,1001,101);
  `device_slave_connections_TB_CONFIG_4(1,1002,102);
  `device_slave_connections_TB_CONFIG_4(1,1003,103);
  `device_slave_connections_TB_CONFIG_4(1,1004,104);
  `device_slave_connections_TB_CONFIG_4(1,1005,105);
  `device_slave_connections_TB_CONFIG_4(1,1006,106);
  `device_slave_connections_TB_CONFIG_4(1,1007,107);
  `device_slave_connections_TB_CONFIG_4(1,1008,108);
  `device_slave_connections_TB_CONFIG_4(1,1009,109);
  `device_slave_connections_TB_CONFIG_4(1,1010,110);
  `device_slave_connections_TB_CONFIG_4(1,1011,111);
  `device_slave_connections_TB_CONFIG_4(1,1012,112);
  `device_slave_connections_TB_CONFIG_4(1,1013,113);
  `device_slave_connections_TB_CONFIG_4(1,1014,114);
  `device_slave_connections_TB_CONFIG_4(1,1015,115);
  `device_slave_connections_TB_CONFIG_4(1,1016,116);
  `device_slave_connections_TB_CONFIG_4(1,1017,117);
  `device_slave_connections_TB_CONFIG_4(1,1018,118);
  `device_slave_connections_TB_CONFIG_4(1,1019,119);
  `device_slave_connections_TB_CONFIG_4(1,1020,120);
  `device_slave_connections_TB_CONFIG_4(1,1021,121);
  `device_slave_connections_TB_CONFIG_4(1,1022,122);
  `device_slave_connections_TB_CONFIG_4(1,1023,123);
  `device_slave_connections_TB_CONFIG_4(1,1024,124);
  `device_slave_connections_TB_CONFIG_4(1,1025,125);
  `device_slave_connections_TB_CONFIG_4(1,1026,126);
  `device_slave_connections_TB_CONFIG_4(1,1027,127);
  `device_slave_connections_TB_CONFIG_4(1,1028,128);
  `device_slave_connections_TB_CONFIG_4(1,1029,129);
  `device_slave_connections_TB_CONFIG_4(1,1030,130);
  `device_slave_connections_TB_CONFIG_4(1,1031,131);
  `device_slave_connections_TB_CONFIG_4(1,1032,132);
  `device_slave_connections_TB_CONFIG_4(1,1033,133);
  `device_slave_connections_TB_CONFIG_4(1,1034,134);
  `device_slave_connections_TB_CONFIG_4(1,1035,135);
  `device_slave_connections_TB_CONFIG_4(1,1036,136);
  `device_slave_connections_TB_CONFIG_4(1,1037,137);
  `device_slave_connections_TB_CONFIG_4(1,1038,138);
  `device_slave_connections_TB_CONFIG_4(1,1039,139);
  `device_slave_connections_TB_CONFIG_4(1,1040,140);
  `device_slave_connections_TB_CONFIG_4(1,1041,141);
  `device_slave_connections_TB_CONFIG_4(1,1042,142);
  `device_slave_connections_TB_CONFIG_4(1,1043,143);
  `device_slave_connections_TB_CONFIG_4(1,1044,144);
  `device_slave_connections_TB_CONFIG_4(1,1045,145);
  `device_slave_connections_TB_CONFIG_4(1,1046,146);
  `device_slave_connections_TB_CONFIG_4(1,1047,147);
  `device_slave_connections_TB_CONFIG_4(1,1048,148);
  `device_slave_connections_TB_CONFIG_4(1,1049,149);
  `device_slave_connections_TB_CONFIG_4(1,1050,150);
  `device_slave_connections_TB_CONFIG_4(1,1051,151);
  `device_slave_connections_TB_CONFIG_4(1,1052,152);
  `device_slave_connections_TB_CONFIG_4(1,1053,153);
  `device_slave_connections_TB_CONFIG_4(1,1054,154);
  `device_slave_connections_TB_CONFIG_4(1,1055,155);
  `device_slave_connections_TB_CONFIG_4(1,1056,156);
  `device_slave_connections_TB_CONFIG_4(1,1057,157);
  `device_slave_connections_TB_CONFIG_4(1,1058,158);
  `device_slave_connections_TB_CONFIG_4(1,1059,159);
  `device_slave_connections_TB_CONFIG_4(1,1060,160);
  `device_slave_connections_TB_CONFIG_4(1,1061,161);
  `device_slave_connections_TB_CONFIG_4(1,1062,162);
  `device_slave_connections_TB_CONFIG_4(1,1063,163);
  `device_slave_connections_TB_CONFIG_4(1,1064,164);
  `device_slave_connections_TB_CONFIG_4(1,1065,165);
  `device_slave_connections_TB_CONFIG_4(1,1066,166);
  `device_slave_connections_TB_CONFIG_4(1,1067,167);
  `device_slave_connections_TB_CONFIG_4(1,1068,168);
  `device_slave_connections_TB_CONFIG_4(1,1069,169);
  `device_slave_connections_TB_CONFIG_4(1,1070,170);
  `device_slave_connections_TB_CONFIG_4(1,1071,171);
  `device_slave_connections_TB_CONFIG_4(1,1072,172);
  `device_slave_connections_TB_CONFIG_4(1,1073,173);
  `device_slave_connections_TB_CONFIG_4(1,1074,174);
  `device_slave_connections_TB_CONFIG_4(1,1075,175);
  `device_slave_connections_TB_CONFIG_4(1,1076,176);
  `device_slave_connections_TB_CONFIG_4(1,1077,177);
  `device_slave_connections_TB_CONFIG_4(1,1078,178);
  `device_slave_connections_TB_CONFIG_4(1,1079,179);
  `device_slave_connections_TB_CONFIG_4(1,1080,180);
  `device_slave_connections_TB_CONFIG_4(1,1081,181);
  `device_slave_connections_TB_CONFIG_4(1,1082,182);
  `device_slave_connections_TB_CONFIG_4(1,1083,183);
  `device_slave_connections_TB_CONFIG_4(1,1084,184);
  `device_slave_connections_TB_CONFIG_4(1,1085,185);
  `device_slave_connections_TB_CONFIG_4(1,1086,186);
  `device_slave_connections_TB_CONFIG_4(1,1087,187);
  `device_slave_connections_TB_CONFIG_4(1,1088,188);
  `device_slave_connections_TB_CONFIG_4(1,1089,189);
  `device_slave_connections_TB_CONFIG_4(1,1090,190);
  `device_slave_connections_TB_CONFIG_4(1,1091,191);
  `device_slave_connections_TB_CONFIG_4(1,1092,192);
  `device_slave_connections_TB_CONFIG_4(1,1093,193);
  `device_slave_connections_TB_CONFIG_4(1,1094,194);
  `device_slave_connections_TB_CONFIG_4(1,1095,195);
  `device_slave_connections_TB_CONFIG_4(1,1096,196);
  `device_slave_connections_TB_CONFIG_4(1,1097,197);
  `device_slave_connections_TB_CONFIG_4(1,1098,198);
  `device_slave_connections_TB_CONFIG_4(1,1099,199);
  `device_slave_connections_TB_CONFIG_4(1,1100,200);
  `device_slave_connections_TB_CONFIG_4(1,1101,201);
  `device_slave_connections_TB_CONFIG_4(1,1102,202);
  `device_slave_connections_TB_CONFIG_4(1,1103,203);
  `device_slave_connections_TB_CONFIG_4(1,1104,204);
  `device_slave_connections_TB_CONFIG_4(1,1105,205);
  `device_slave_connections_TB_CONFIG_4(1,1106,206);
  `device_slave_connections_TB_CONFIG_4(1,1107,207);
  `device_slave_connections_TB_CONFIG_4(1,1108,208);
  `device_slave_connections_TB_CONFIG_4(1,1109,209);
  `device_slave_connections_TB_CONFIG_4(1,1110,210);
  `device_slave_connections_TB_CONFIG_4(1,1111,211);
  `device_slave_connections_TB_CONFIG_4(1,1112,212);
  `device_slave_connections_TB_CONFIG_4(1,1113,213);
  `device_slave_connections_TB_CONFIG_4(1,1114,214);
  `device_slave_connections_TB_CONFIG_4(1,1115,215);
  `device_slave_connections_TB_CONFIG_4(1,1116,216);
  `device_slave_connections_TB_CONFIG_4(1,1117,217);
  `device_slave_connections_TB_CONFIG_4(1,1118,218);
  `device_slave_connections_TB_CONFIG_4(1,1119,219);
  `device_slave_connections_TB_CONFIG_4(1,1120,220);
  `device_slave_connections_TB_CONFIG_4(1,1121,221);
  `device_slave_connections_TB_CONFIG_4(1,1122,222);
  `device_slave_connections_TB_CONFIG_4(1,1123,223);
  `device_slave_connections_TB_CONFIG_4(1,1124,224);
  `device_slave_connections_TB_CONFIG_4(1,1125,225);
  `device_slave_connections_TB_CONFIG_4(1,1126,226);
  `device_slave_connections_TB_CONFIG_4(1,1127,227);
  `device_slave_connections_TB_CONFIG_4(1,1128,228);
  `device_slave_connections_TB_CONFIG_4(1,1129,229);
  `device_slave_connections_TB_CONFIG_4(1,1130,230);
  `device_slave_connections_TB_CONFIG_4(1,1131,231);
  `device_slave_connections_TB_CONFIG_4(1,1132,232);
  `device_slave_connections_TB_CONFIG_4(1,1133,233);
  `device_slave_connections_TB_CONFIG_4(1,1134,234);
  `device_slave_connections_TB_CONFIG_4(1,1135,235);
  `device_slave_connections_TB_CONFIG_4(1,1136,236);
  `device_slave_connections_TB_CONFIG_4(1,1137,237);
  `device_slave_connections_TB_CONFIG_4(1,1138,238);
  `device_slave_connections_TB_CONFIG_4(1,1139,239);
  `device_slave_connections_TB_CONFIG_4(1,1140,240);
  `device_slave_connections_TB_CONFIG_4(1,1141,241);
  `device_slave_connections_TB_CONFIG_4(1,1142,242);
  `device_slave_connections_TB_CONFIG_4(1,1143,243);
  `device_slave_connections_TB_CONFIG_4(1,1144,244);
  `device_slave_connections_TB_CONFIG_4(1,1145,245);
  `device_slave_connections_TB_CONFIG_4(1,1146,246);
  `device_slave_connections_TB_CONFIG_4(1,1147,247);
  `device_slave_connections_TB_CONFIG_4(1,1148,248);
  `device_slave_connections_TB_CONFIG_4(1,1149,249);
  `device_slave_connections_TB_CONFIG_4(1,1150,250);
  `device_slave_connections_TB_CONFIG_4(1,1151,251);
  `device_slave_connections_TB_CONFIG_4(1,1152,252);
  `device_slave_connections_TB_CONFIG_4(1,1153,253);
  `device_slave_connections_TB_CONFIG_4(1,1154,254);
  `device_slave_connections_TB_CONFIG_4(1,1155,255);
  `device_slave_connections_TB_CONFIG_4(1,1156,256);
  `device_slave_connections_TB_CONFIG_4(1,1157,257);
  `device_slave_connections_TB_CONFIG_4(1,1158,258);
  `device_slave_connections_TB_CONFIG_4(1,1159,259);
  `device_slave_connections_TB_CONFIG_4(1,1160,260);
  `device_slave_connections_TB_CONFIG_4(1,1161,261);
  `device_slave_connections_TB_CONFIG_4(1,1162,262);
  `device_slave_connections_TB_CONFIG_4(1,1163,263);
  `device_slave_connections_TB_CONFIG_4(1,1164,264);
  `device_slave_connections_TB_CONFIG_4(1,1165,265);
  `device_slave_connections_TB_CONFIG_4(1,1166,266);
  `device_slave_connections_TB_CONFIG_4(1,1167,267);
  `device_slave_connections_TB_CONFIG_4(1,1168,268);
  `device_slave_connections_TB_CONFIG_4(1,1169,269);
  `device_slave_connections_TB_CONFIG_4(1,1170,270);
  `device_slave_connections_TB_CONFIG_4(1,1171,271);
  `device_slave_connections_TB_CONFIG_4(1,1172,272);
  `device_slave_connections_TB_CONFIG_4(1,1173,273);
  `device_slave_connections_TB_CONFIG_4(1,1174,274);
  `device_slave_connections_TB_CONFIG_4(1,1175,275);
  `device_slave_connections_TB_CONFIG_4(1,1176,276);
  `device_slave_connections_TB_CONFIG_4(1,1177,277);
  `device_slave_connections_TB_CONFIG_4(1,1178,278);
  `device_slave_connections_TB_CONFIG_4(1,1179,279);
  `device_slave_connections_TB_CONFIG_4(1,1180,280);
  `device_slave_connections_TB_CONFIG_4(1,1181,281);
  `device_slave_connections_TB_CONFIG_4(1,1182,282);
  `device_slave_connections_TB_CONFIG_4(1,1183,283);
  `device_slave_connections_TB_CONFIG_4(1,1184,284);
  `device_slave_connections_TB_CONFIG_4(1,1185,285);
  `device_slave_connections_TB_CONFIG_4(1,1186,286);
  `device_slave_connections_TB_CONFIG_4(1,1187,287);
  `device_slave_connections_TB_CONFIG_4(1,1188,288);
  `device_slave_connections_TB_CONFIG_4(1,1189,289);
  `device_slave_connections_TB_CONFIG_4(1,1190,290);
  `device_slave_connections_TB_CONFIG_4(1,1191,291);
  `device_slave_connections_TB_CONFIG_4(1,1192,292);
  `device_slave_connections_TB_CONFIG_4(1,1193,293);
  `device_slave_connections_TB_CONFIG_4(1,1194,294);
  `device_slave_connections_TB_CONFIG_4(1,1195,295);
  `device_slave_connections_TB_CONFIG_4(1,1196,296);
  `device_slave_connections_TB_CONFIG_4(1,1197,297);
  `device_slave_connections_TB_CONFIG_4(1,1198,298);
  `device_slave_connections_TB_CONFIG_4(1,1199,299);
  `device_slave_connections_TB_CONFIG_4(1,1200,300);
  `device_slave_connections_TB_CONFIG_4(1,1201,301);
  `device_slave_connections_TB_CONFIG_4(1,1202,302);
  `device_slave_connections_TB_CONFIG_4(1,1203,303);
  `device_slave_connections_TB_CONFIG_4(1,1204,304);
  `device_slave_connections_TB_CONFIG_4(1,1205,305);
  `device_slave_connections_TB_CONFIG_4(1,1206,306);
  `device_slave_connections_TB_CONFIG_4(1,1207,307);
  `device_slave_connections_TB_CONFIG_4(1,1208,308);
  `device_slave_connections_TB_CONFIG_4(1,1209,309);
  `device_slave_connections_TB_CONFIG_4(1,1210,310);
  `device_slave_connections_TB_CONFIG_4(1,1211,311);
  `device_slave_connections_TB_CONFIG_4(1,1212,312);
  `device_slave_connections_TB_CONFIG_4(1,1213,313);
  `device_slave_connections_TB_CONFIG_4(1,1214,314);
  `device_slave_connections_TB_CONFIG_4(1,1215,315);
  `device_slave_connections_TB_CONFIG_4(1,1216,316);
  `device_slave_connections_TB_CONFIG_4(1,1217,317);
  `device_slave_connections_TB_CONFIG_4(1,1218,318);
  `device_slave_connections_TB_CONFIG_4(1,1219,319);
  `device_slave_connections_TB_CONFIG_4(1,1220,320);
  `device_slave_connections_TB_CONFIG_4(1,1221,321);
  `device_slave_connections_TB_CONFIG_4(1,1222,322);
  `device_slave_connections_TB_CONFIG_4(1,1223,323);
  `device_slave_connections_TB_CONFIG_4(1,1224,324);
  `device_slave_connections_TB_CONFIG_4(1,1225,325);
  `device_slave_connections_TB_CONFIG_4(1,1226,326);
  `device_slave_connections_TB_CONFIG_4(1,1227,327);
  `device_slave_connections_TB_CONFIG_4(1,1228,328);
  `device_slave_connections_TB_CONFIG_4(1,1229,329);
  `device_slave_connections_TB_CONFIG_4(1,1230,330);
  `device_slave_connections_TB_CONFIG_4(1,1231,331);
  `device_slave_connections_TB_CONFIG_4(1,1232,332);
  `device_slave_connections_TB_CONFIG_4(1,1233,333);
  `device_slave_connections_TB_CONFIG_4(1,1234,334);
  `device_slave_connections_TB_CONFIG_4(1,1235,335);
  `device_slave_connections_TB_CONFIG_4(1,1236,336);
  `device_slave_connections_TB_CONFIG_4(1,1237,337);
  `device_slave_connections_TB_CONFIG_4(1,1238,338);
  `device_slave_connections_TB_CONFIG_4(1,1239,339);
  `device_slave_connections_TB_CONFIG_4(1,1240,340);
  `device_slave_connections_TB_CONFIG_4(1,1241,341);
  `device_slave_connections_TB_CONFIG_4(1,1242,342);
  `device_slave_connections_TB_CONFIG_4(1,1243,343);
  `device_slave_connections_TB_CONFIG_4(1,1244,344);
  `device_slave_connections_TB_CONFIG_4(1,1245,345);
  `device_slave_connections_TB_CONFIG_4(1,1246,346);
  `device_slave_connections_TB_CONFIG_4(1,1247,347);
  `device_slave_connections_TB_CONFIG_4(1,1248,348);
  `device_slave_connections_TB_CONFIG_4(1,1249,349);
  `device_slave_connections_TB_CONFIG_4(1,1250,350);
  `device_slave_connections_TB_CONFIG_4(1,1251,351);
  `device_slave_connections_TB_CONFIG_4(1,1252,352);
  `device_slave_connections_TB_CONFIG_4(1,1253,353);
  `device_slave_connections_TB_CONFIG_4(1,1254,354);
  `device_slave_connections_TB_CONFIG_4(1,1255,355);
  `device_slave_connections_TB_CONFIG_4(1,1256,356);
  `device_slave_connections_TB_CONFIG_4(1,1257,357);
  `device_slave_connections_TB_CONFIG_4(1,1258,358);
  `device_slave_connections_TB_CONFIG_4(1,1259,359);
  `device_slave_connections_TB_CONFIG_4(1,1260,360);
  `device_slave_connections_TB_CONFIG_4(1,1261,361);
  `device_slave_connections_TB_CONFIG_4(1,1262,362);
  `device_slave_connections_TB_CONFIG_4(1,1263,363);
  `device_slave_connections_TB_CONFIG_4(1,1264,364);
  `device_slave_connections_TB_CONFIG_4(1,1265,365);
  `device_slave_connections_TB_CONFIG_4(1,1266,366);
  `device_slave_connections_TB_CONFIG_4(1,1267,367);
  `device_slave_connections_TB_CONFIG_4(1,1268,368);
  `device_slave_connections_TB_CONFIG_4(1,1269,369);
  `device_slave_connections_TB_CONFIG_4(1,1270,370);
  `device_slave_connections_TB_CONFIG_4(1,1271,371);
  `device_slave_connections_TB_CONFIG_4(1,1272,372);
  `device_slave_connections_TB_CONFIG_4(1,1273,373);
  `device_slave_connections_TB_CONFIG_4(1,1274,374);
  `device_slave_connections_TB_CONFIG_4(1,1275,375);
  `device_slave_connections_TB_CONFIG_4(1,1276,376);
  `device_slave_connections_TB_CONFIG_4(1,1277,377);
  `device_slave_connections_TB_CONFIG_4(1,1278,378);
  `device_slave_connections_TB_CONFIG_4(1,1279,379);
  `device_slave_connections_TB_CONFIG_4(1,1280,380);
  `device_slave_connections_TB_CONFIG_4(1,1281,381);
  `device_slave_connections_TB_CONFIG_4(1,1282,382);
  `device_slave_connections_TB_CONFIG_4(1,1283,383);
  `device_slave_connections_TB_CONFIG_4(1,1284,384);
  `device_slave_connections_TB_CONFIG_4(1,1285,385);
  `device_slave_connections_TB_CONFIG_4(1,1286,386);
  `device_slave_connections_TB_CONFIG_4(1,1287,387);
  `device_slave_connections_TB_CONFIG_4(1,1288,388);
  `device_slave_connections_TB_CONFIG_4(1,1289,389);
  `device_slave_connections_TB_CONFIG_4(1,1290,390);
  `device_slave_connections_TB_CONFIG_4(1,1291,391);
  `device_slave_connections_TB_CONFIG_4(1,1292,392);
  `device_slave_connections_TB_CONFIG_4(1,1293,393);
  `device_slave_connections_TB_CONFIG_4(1,1294,394);
  `device_slave_connections_TB_CONFIG_4(1,1295,395);
  `device_slave_connections_TB_CONFIG_4(1,1296,396);
  `device_slave_connections_TB_CONFIG_4(1,1297,397);
  `device_slave_connections_TB_CONFIG_4(1,1298,398);
  `device_slave_connections_TB_CONFIG_4(1,1299,399);
  `device_slave_connections_TB_CONFIG_4(1,1300,400);
  `device_slave_connections_TB_CONFIG_4(1,1301,401);
  `device_slave_connections_TB_CONFIG_4(1,1302,402);
  `device_slave_connections_TB_CONFIG_4(1,1303,403);
  `device_slave_connections_TB_CONFIG_4(1,1304,404);
  `device_slave_connections_TB_CONFIG_4(1,1305,405);
  `device_slave_connections_TB_CONFIG_4(1,1306,406);
  `device_slave_connections_TB_CONFIG_4(1,1307,407);
  `device_slave_connections_TB_CONFIG_4(1,1308,408);
  `device_slave_connections_TB_CONFIG_4(1,1309,409);
  `device_slave_connections_TB_CONFIG_4(1,1310,410);
  `device_slave_connections_TB_CONFIG_4(1,1311,411);
  `device_slave_connections_TB_CONFIG_4(1,1312,412);
  `device_slave_connections_TB_CONFIG_4(1,1313,413);
  `device_slave_connections_TB_CONFIG_4(1,1314,414);
  `device_slave_connections_TB_CONFIG_4(1,1315,415);
  `device_slave_connections_TB_CONFIG_4(1,1316,416);
  `device_slave_connections_TB_CONFIG_4(1,1317,417);
  `device_slave_connections_TB_CONFIG_4(1,1318,418);
  `device_slave_connections_TB_CONFIG_4(1,1319,419);
  `device_slave_connections_TB_CONFIG_4(1,1320,420);
  `device_slave_connections_TB_CONFIG_4(1,1321,421);
  `device_slave_connections_TB_CONFIG_4(1,1322,422);
  `device_slave_connections_TB_CONFIG_4(1,1323,423);
  `device_slave_connections_TB_CONFIG_4(1,1324,424);
  `device_slave_connections_TB_CONFIG_4(1,1325,425);
  `device_slave_connections_TB_CONFIG_4(1,1326,426);
  `device_slave_connections_TB_CONFIG_4(1,1327,427);
  `device_slave_connections_TB_CONFIG_4(1,1328,428);
  `device_slave_connections_TB_CONFIG_4(1,1329,429);
  `device_slave_connections_TB_CONFIG_4(1,1330,430);
  `device_slave_connections_TB_CONFIG_4(1,1331,431);
  `device_slave_connections_TB_CONFIG_4(1,1332,432);
  `device_slave_connections_TB_CONFIG_4(1,1333,433);
  `device_slave_connections_TB_CONFIG_4(1,1334,434);
  `device_slave_connections_TB_CONFIG_4(1,1335,435);
  `device_slave_connections_TB_CONFIG_4(1,1336,436);
  `device_slave_connections_TB_CONFIG_4(1,1337,437);
  `device_slave_connections_TB_CONFIG_4(1,1338,438);
  `device_slave_connections_TB_CONFIG_4(1,1339,439);
  `device_slave_connections_TB_CONFIG_4(1,1340,440);
  `device_slave_connections_TB_CONFIG_4(1,1341,441);
  `device_slave_connections_TB_CONFIG_4(1,1342,442);
  `device_slave_connections_TB_CONFIG_4(1,1343,443);
  `device_slave_connections_TB_CONFIG_4(1,1344,444);
  `device_slave_connections_TB_CONFIG_4(1,1345,445);
  `device_slave_connections_TB_CONFIG_4(1,1346,446);
  `device_slave_connections_TB_CONFIG_4(1,1347,447);
  `device_slave_connections_TB_CONFIG_4(1,1348,448);
  `device_slave_connections_TB_CONFIG_4(1,1349,449);
	`device_slave_connections_TB_CONFIG_4(2,1350,0);
  `device_slave_connections_TB_CONFIG_4(2,1351,1);
  `device_slave_connections_TB_CONFIG_4(2,1352,2);
  `device_slave_connections_TB_CONFIG_4(2,1353,3);
  `device_slave_connections_TB_CONFIG_4(2,1354,4);
  `device_slave_connections_TB_CONFIG_4(2,1355,5);
  `device_slave_connections_TB_CONFIG_4(2,1356,6);
  `device_slave_connections_TB_CONFIG_4(2,1357,7);
  `device_slave_connections_TB_CONFIG_4(2,1358,8);
  `device_slave_connections_TB_CONFIG_4(2,1359,9);
  `device_slave_connections_TB_CONFIG_4(2,1360,10);
  `device_slave_connections_TB_CONFIG_4(2,1361,11);
  `device_slave_connections_TB_CONFIG_4(2,1362,12);
  `device_slave_connections_TB_CONFIG_4(2,1363,13);
  `device_slave_connections_TB_CONFIG_4(2,1364,14);
  `device_slave_connections_TB_CONFIG_4(2,1365,15);
  `device_slave_connections_TB_CONFIG_4(2,1366,16);
  `device_slave_connections_TB_CONFIG_4(2,1367,17);
  `device_slave_connections_TB_CONFIG_4(2,1368,18);
  `device_slave_connections_TB_CONFIG_4(2,1369,19);
  `device_slave_connections_TB_CONFIG_4(2,1370,20);
  `device_slave_connections_TB_CONFIG_4(2,1371,21);
  `device_slave_connections_TB_CONFIG_4(2,1372,22);
  `device_slave_connections_TB_CONFIG_4(2,1373,23);
  `device_slave_connections_TB_CONFIG_4(2,1374,24);
  `device_slave_connections_TB_CONFIG_4(2,1375,25);
  `device_slave_connections_TB_CONFIG_4(2,1376,26);
  `device_slave_connections_TB_CONFIG_4(2,1377,27);
  `device_slave_connections_TB_CONFIG_4(2,1378,28);
  `device_slave_connections_TB_CONFIG_4(2,1379,29);
  `device_slave_connections_TB_CONFIG_4(2,1380,30);
  `device_slave_connections_TB_CONFIG_4(2,1381,31);
  `device_slave_connections_TB_CONFIG_4(2,1382,32);
  `device_slave_connections_TB_CONFIG_4(2,1383,33);
  `device_slave_connections_TB_CONFIG_4(2,1384,34);
  `device_slave_connections_TB_CONFIG_4(2,1385,35);
  `device_slave_connections_TB_CONFIG_4(2,1386,36);
  `device_slave_connections_TB_CONFIG_4(2,1387,37);
  `device_slave_connections_TB_CONFIG_4(2,1388,38);
  `device_slave_connections_TB_CONFIG_4(2,1389,39);
  `device_slave_connections_TB_CONFIG_4(2,1390,40);
  `device_slave_connections_TB_CONFIG_4(2,1391,41);
  `device_slave_connections_TB_CONFIG_4(2,1392,42);
  `device_slave_connections_TB_CONFIG_4(2,1393,43);
  `device_slave_connections_TB_CONFIG_4(2,1394,44);
  `device_slave_connections_TB_CONFIG_4(2,1395,45);
  `device_slave_connections_TB_CONFIG_4(2,1396,46);
  `device_slave_connections_TB_CONFIG_4(2,1397,47);
  `device_slave_connections_TB_CONFIG_4(2,1398,48);
  `device_slave_connections_TB_CONFIG_4(2,1399,49);
  `device_slave_connections_TB_CONFIG_4(2,1400,50);
  `device_slave_connections_TB_CONFIG_4(2,1401,51);
  `device_slave_connections_TB_CONFIG_4(2,1402,52);
  `device_slave_connections_TB_CONFIG_4(2,1403,53);
  `device_slave_connections_TB_CONFIG_4(2,1404,54);
  `device_slave_connections_TB_CONFIG_4(2,1405,55);
  `device_slave_connections_TB_CONFIG_4(2,1406,56);
  `device_slave_connections_TB_CONFIG_4(2,1407,57);
  `device_slave_connections_TB_CONFIG_4(2,1408,58);
  `device_slave_connections_TB_CONFIG_4(2,1409,59);
  `device_slave_connections_TB_CONFIG_4(2,1410,60);
  `device_slave_connections_TB_CONFIG_4(2,1411,61);
  `device_slave_connections_TB_CONFIG_4(2,1412,62);
  `device_slave_connections_TB_CONFIG_4(2,1413,63);
  `device_slave_connections_TB_CONFIG_4(2,1414,64);
  `device_slave_connections_TB_CONFIG_4(2,1415,65);
  `device_slave_connections_TB_CONFIG_4(2,1416,66);
  `device_slave_connections_TB_CONFIG_4(2,1417,67);
  `device_slave_connections_TB_CONFIG_4(2,1418,68);
  `device_slave_connections_TB_CONFIG_4(2,1419,69);
  `device_slave_connections_TB_CONFIG_4(2,1420,70);
  `device_slave_connections_TB_CONFIG_4(2,1421,71);
  `device_slave_connections_TB_CONFIG_4(2,1422,72);
  `device_slave_connections_TB_CONFIG_4(2,1423,73);
  `device_slave_connections_TB_CONFIG_4(2,1424,74);
  `device_slave_connections_TB_CONFIG_4(2,1425,75);
  `device_slave_connections_TB_CONFIG_4(2,1426,76);
  `device_slave_connections_TB_CONFIG_4(2,1427,77);
  `device_slave_connections_TB_CONFIG_4(2,1428,78);
  `device_slave_connections_TB_CONFIG_4(2,1429,79);
  `device_slave_connections_TB_CONFIG_4(2,1430,80);
  `device_slave_connections_TB_CONFIG_4(2,1431,81);
  `device_slave_connections_TB_CONFIG_4(2,1432,82);
  `device_slave_connections_TB_CONFIG_4(2,1433,83);
  `device_slave_connections_TB_CONFIG_4(2,1434,84);
  `device_slave_connections_TB_CONFIG_4(2,1435,85);
  `device_slave_connections_TB_CONFIG_4(2,1436,86);
  `device_slave_connections_TB_CONFIG_4(2,1437,87);
  `device_slave_connections_TB_CONFIG_4(2,1438,88);
  `device_slave_connections_TB_CONFIG_4(2,1439,89);
  `device_slave_connections_TB_CONFIG_4(2,1440,90);
  `device_slave_connections_TB_CONFIG_4(2,1441,91);
  `device_slave_connections_TB_CONFIG_4(2,1442,92);
  `device_slave_connections_TB_CONFIG_4(2,1443,93);
  `device_slave_connections_TB_CONFIG_4(2,1444,94);
  `device_slave_connections_TB_CONFIG_4(2,1445,95);
  `device_slave_connections_TB_CONFIG_4(2,1446,96);
  `device_slave_connections_TB_CONFIG_4(2,1447,97);
  `device_slave_connections_TB_CONFIG_4(2,1448,98);
  `device_slave_connections_TB_CONFIG_4(2,1449,99);
  `device_slave_connections_TB_CONFIG_4(2,1450,100);
  `device_slave_connections_TB_CONFIG_4(2,1451,101);
  `device_slave_connections_TB_CONFIG_4(2,1452,102);
  `device_slave_connections_TB_CONFIG_4(2,1453,103);
  `device_slave_connections_TB_CONFIG_4(2,1454,104);
  `device_slave_connections_TB_CONFIG_4(2,1455,105);
  `device_slave_connections_TB_CONFIG_4(2,1456,106);
  `device_slave_connections_TB_CONFIG_4(2,1457,107);
  `device_slave_connections_TB_CONFIG_4(2,1458,108);
  `device_slave_connections_TB_CONFIG_4(2,1459,109);
  `device_slave_connections_TB_CONFIG_4(2,1460,110);
  `device_slave_connections_TB_CONFIG_4(2,1461,111);
  `device_slave_connections_TB_CONFIG_4(2,1462,112);
  `device_slave_connections_TB_CONFIG_4(2,1463,113);
  `device_slave_connections_TB_CONFIG_4(2,1464,114);
  `device_slave_connections_TB_CONFIG_4(2,1465,115);
  `device_slave_connections_TB_CONFIG_4(2,1466,116);
  `device_slave_connections_TB_CONFIG_4(2,1467,117);
  `device_slave_connections_TB_CONFIG_4(2,1468,118);
  `device_slave_connections_TB_CONFIG_4(2,1469,119);
  `device_slave_connections_TB_CONFIG_4(2,1470,120);
  `device_slave_connections_TB_CONFIG_4(2,1471,121);
  `device_slave_connections_TB_CONFIG_4(2,1472,122);
  `device_slave_connections_TB_CONFIG_4(2,1473,123);
  `device_slave_connections_TB_CONFIG_4(2,1474,124);
  `device_slave_connections_TB_CONFIG_4(2,1475,125);
  `device_slave_connections_TB_CONFIG_4(2,1476,126);
  `device_slave_connections_TB_CONFIG_4(2,1477,127);
  `device_slave_connections_TB_CONFIG_4(2,1478,128);
  `device_slave_connections_TB_CONFIG_4(2,1479,129);
  `device_slave_connections_TB_CONFIG_4(2,1480,130);
  `device_slave_connections_TB_CONFIG_4(2,1481,131);
  `device_slave_connections_TB_CONFIG_4(2,1482,132);
  `device_slave_connections_TB_CONFIG_4(2,1483,133);
  `device_slave_connections_TB_CONFIG_4(2,1484,134);
  `device_slave_connections_TB_CONFIG_4(2,1485,135);
  `device_slave_connections_TB_CONFIG_4(2,1486,136);
  `device_slave_connections_TB_CONFIG_4(2,1487,137);
  `device_slave_connections_TB_CONFIG_4(2,1488,138);
  `device_slave_connections_TB_CONFIG_4(2,1489,139);
  `device_slave_connections_TB_CONFIG_4(2,1490,140);
  `device_slave_connections_TB_CONFIG_4(2,1491,141);
  `device_slave_connections_TB_CONFIG_4(2,1492,142);
  `device_slave_connections_TB_CONFIG_4(2,1493,143);
  `device_slave_connections_TB_CONFIG_4(2,1494,144);
  `device_slave_connections_TB_CONFIG_4(2,1495,145);
  `device_slave_connections_TB_CONFIG_4(2,1496,146);
  `device_slave_connections_TB_CONFIG_4(2,1497,147);
  `device_slave_connections_TB_CONFIG_4(2,1498,148);
  `device_slave_connections_TB_CONFIG_4(2,1499,149);
  `device_slave_connections_TB_CONFIG_4(2,1500,150);
  `device_slave_connections_TB_CONFIG_4(2,1501,151);
  `device_slave_connections_TB_CONFIG_4(2,1502,152);
  `device_slave_connections_TB_CONFIG_4(2,1503,153);
  `device_slave_connections_TB_CONFIG_4(2,1504,154);
  `device_slave_connections_TB_CONFIG_4(2,1505,155);
  `device_slave_connections_TB_CONFIG_4(2,1506,156);
  `device_slave_connections_TB_CONFIG_4(2,1507,157);
  `device_slave_connections_TB_CONFIG_4(2,1508,158);
  `device_slave_connections_TB_CONFIG_4(2,1509,159);
  `device_slave_connections_TB_CONFIG_4(2,1510,160);
  `device_slave_connections_TB_CONFIG_4(2,1511,161);
  `device_slave_connections_TB_CONFIG_4(2,1512,162);
  `device_slave_connections_TB_CONFIG_4(2,1513,163);
  `device_slave_connections_TB_CONFIG_4(2,1514,164);
  `device_slave_connections_TB_CONFIG_4(2,1515,165);
  `device_slave_connections_TB_CONFIG_4(2,1516,166);
  `device_slave_connections_TB_CONFIG_4(2,1517,167);
  `device_slave_connections_TB_CONFIG_4(2,1518,168);
  `device_slave_connections_TB_CONFIG_4(2,1519,169);
  `device_slave_connections_TB_CONFIG_4(2,1520,170);
  `device_slave_connections_TB_CONFIG_4(2,1521,171);
  `device_slave_connections_TB_CONFIG_4(2,1522,172);
  `device_slave_connections_TB_CONFIG_4(2,1523,173);
  `device_slave_connections_TB_CONFIG_4(2,1524,174);
  `device_slave_connections_TB_CONFIG_4(2,1525,175);
  `device_slave_connections_TB_CONFIG_4(2,1526,176);
  `device_slave_connections_TB_CONFIG_4(2,1527,177);
  `device_slave_connections_TB_CONFIG_4(2,1528,178);
  `device_slave_connections_TB_CONFIG_4(2,1529,179);
  `device_slave_connections_TB_CONFIG_4(2,1530,180);
  `device_slave_connections_TB_CONFIG_4(2,1531,181);
  `device_slave_connections_TB_CONFIG_4(2,1532,182);
  `device_slave_connections_TB_CONFIG_4(2,1533,183);
  `device_slave_connections_TB_CONFIG_4(2,1534,184);
  `device_slave_connections_TB_CONFIG_4(2,1535,185);
  `device_slave_connections_TB_CONFIG_4(2,1536,186);
  `device_slave_connections_TB_CONFIG_4(2,1537,187);
  `device_slave_connections_TB_CONFIG_4(2,1538,188);
  `device_slave_connections_TB_CONFIG_4(2,1539,189);
  `device_slave_connections_TB_CONFIG_4(2,1540,190);
  `device_slave_connections_TB_CONFIG_4(2,1541,191);
  `device_slave_connections_TB_CONFIG_4(2,1542,192);
  `device_slave_connections_TB_CONFIG_4(2,1543,193);
  `device_slave_connections_TB_CONFIG_4(2,1544,194);
  `device_slave_connections_TB_CONFIG_4(2,1545,195);
  `device_slave_connections_TB_CONFIG_4(2,1546,196);
  `device_slave_connections_TB_CONFIG_4(2,1547,197);
  `device_slave_connections_TB_CONFIG_4(2,1548,198);
  `device_slave_connections_TB_CONFIG_4(2,1549,199);
  `device_slave_connections_TB_CONFIG_4(2,1550,200);
  `device_slave_connections_TB_CONFIG_4(2,1551,201);
  `device_slave_connections_TB_CONFIG_4(2,1552,202);
  `device_slave_connections_TB_CONFIG_4(2,1553,203);
  `device_slave_connections_TB_CONFIG_4(2,1554,204);
  `device_slave_connections_TB_CONFIG_4(2,1555,205);
  `device_slave_connections_TB_CONFIG_4(2,1556,206);
  `device_slave_connections_TB_CONFIG_4(2,1557,207);
  `device_slave_connections_TB_CONFIG_4(2,1558,208);
  `device_slave_connections_TB_CONFIG_4(2,1559,209);
  `device_slave_connections_TB_CONFIG_4(2,1560,210);
  `device_slave_connections_TB_CONFIG_4(2,1561,211);
  `device_slave_connections_TB_CONFIG_4(2,1562,212);
  `device_slave_connections_TB_CONFIG_4(2,1563,213);
  `device_slave_connections_TB_CONFIG_4(2,1564,214);
  `device_slave_connections_TB_CONFIG_4(2,1565,215);
  `device_slave_connections_TB_CONFIG_4(2,1566,216);
  `device_slave_connections_TB_CONFIG_4(2,1567,217);
  `device_slave_connections_TB_CONFIG_4(2,1568,218);
  `device_slave_connections_TB_CONFIG_4(2,1569,219);
  `device_slave_connections_TB_CONFIG_4(2,1570,220);
  `device_slave_connections_TB_CONFIG_4(2,1571,221);
  `device_slave_connections_TB_CONFIG_4(2,1572,222);
  `device_slave_connections_TB_CONFIG_4(2,1573,223);
  `device_slave_connections_TB_CONFIG_4(2,1574,224);
  `device_slave_connections_TB_CONFIG_4(2,1575,225);
  `device_slave_connections_TB_CONFIG_4(2,1576,226);
  `device_slave_connections_TB_CONFIG_4(2,1577,227);
  `device_slave_connections_TB_CONFIG_4(2,1578,228);
  `device_slave_connections_TB_CONFIG_4(2,1579,229);
  `device_slave_connections_TB_CONFIG_4(2,1580,230);
  `device_slave_connections_TB_CONFIG_4(2,1581,231);
  `device_slave_connections_TB_CONFIG_4(2,1582,232);
  `device_slave_connections_TB_CONFIG_4(2,1583,233);
  `device_slave_connections_TB_CONFIG_4(2,1584,234);
  `device_slave_connections_TB_CONFIG_4(2,1585,235);
  `device_slave_connections_TB_CONFIG_4(2,1586,236);
  `device_slave_connections_TB_CONFIG_4(2,1587,237);
  `device_slave_connections_TB_CONFIG_4(2,1588,238);
  `device_slave_connections_TB_CONFIG_4(2,1589,239);
  `device_slave_connections_TB_CONFIG_4(2,1590,240);
  `device_slave_connections_TB_CONFIG_4(2,1591,241);
  `device_slave_connections_TB_CONFIG_4(2,1592,242);
  `device_slave_connections_TB_CONFIG_4(2,1593,243);
  `device_slave_connections_TB_CONFIG_4(2,1594,244);
  `device_slave_connections_TB_CONFIG_4(2,1595,245);
  `device_slave_connections_TB_CONFIG_4(2,1596,246);
  `device_slave_connections_TB_CONFIG_4(2,1597,247);
  `device_slave_connections_TB_CONFIG_4(2,1598,248);
  `device_slave_connections_TB_CONFIG_4(2,1599,249);
  `device_slave_connections_TB_CONFIG_4(2,1600,250);
  `device_slave_connections_TB_CONFIG_4(2,1601,251);
  `device_slave_connections_TB_CONFIG_4(2,1602,252);
  `device_slave_connections_TB_CONFIG_4(2,1603,253);
  `device_slave_connections_TB_CONFIG_4(2,1604,254);
  `device_slave_connections_TB_CONFIG_4(2,1605,255);
  `device_slave_connections_TB_CONFIG_4(2,1606,256);
  `device_slave_connections_TB_CONFIG_4(2,1607,257);
  `device_slave_connections_TB_CONFIG_4(2,1608,258);
  `device_slave_connections_TB_CONFIG_4(2,1609,259);
  `device_slave_connections_TB_CONFIG_4(2,1610,260);
  `device_slave_connections_TB_CONFIG_4(2,1611,261);
  `device_slave_connections_TB_CONFIG_4(2,1612,262);
  `device_slave_connections_TB_CONFIG_4(2,1613,263);
  `device_slave_connections_TB_CONFIG_4(2,1614,264);
  `device_slave_connections_TB_CONFIG_4(2,1615,265);
  `device_slave_connections_TB_CONFIG_4(2,1616,266);
  `device_slave_connections_TB_CONFIG_4(2,1617,267);
  `device_slave_connections_TB_CONFIG_4(2,1618,268);
  `device_slave_connections_TB_CONFIG_4(2,1619,269);
  `device_slave_connections_TB_CONFIG_4(2,1620,270);
  `device_slave_connections_TB_CONFIG_4(2,1621,271);
  `device_slave_connections_TB_CONFIG_4(2,1622,272);
  `device_slave_connections_TB_CONFIG_4(2,1623,273);
  `device_slave_connections_TB_CONFIG_4(2,1624,274);
  `device_slave_connections_TB_CONFIG_4(2,1625,275);
  `device_slave_connections_TB_CONFIG_4(2,1626,276);
  `device_slave_connections_TB_CONFIG_4(2,1627,277);
  `device_slave_connections_TB_CONFIG_4(2,1628,278);
  `device_slave_connections_TB_CONFIG_4(2,1629,279);
  `device_slave_connections_TB_CONFIG_4(2,1630,280);
  `device_slave_connections_TB_CONFIG_4(2,1631,281);
  `device_slave_connections_TB_CONFIG_4(2,1632,282);
  `device_slave_connections_TB_CONFIG_4(2,1633,283);
  `device_slave_connections_TB_CONFIG_4(2,1634,284);
  `device_slave_connections_TB_CONFIG_4(2,1635,285);
  `device_slave_connections_TB_CONFIG_4(2,1636,286);
  `device_slave_connections_TB_CONFIG_4(2,1637,287);
  `device_slave_connections_TB_CONFIG_4(2,1638,288);
  `device_slave_connections_TB_CONFIG_4(2,1639,289);
  `device_slave_connections_TB_CONFIG_4(2,1640,290);
  `device_slave_connections_TB_CONFIG_4(2,1641,291);
  `device_slave_connections_TB_CONFIG_4(2,1642,292);
  `device_slave_connections_TB_CONFIG_4(2,1643,293);
  `device_slave_connections_TB_CONFIG_4(2,1644,294);
  `device_slave_connections_TB_CONFIG_4(2,1645,295);
  `device_slave_connections_TB_CONFIG_4(2,1646,296);
  `device_slave_connections_TB_CONFIG_4(2,1647,297);
  `device_slave_connections_TB_CONFIG_4(2,1648,298);
  `device_slave_connections_TB_CONFIG_4(2,1649,299);
  `device_slave_connections_TB_CONFIG_4(2,1650,300);
  `device_slave_connections_TB_CONFIG_4(2,1651,301);
  `device_slave_connections_TB_CONFIG_4(2,1652,302);
  `device_slave_connections_TB_CONFIG_4(2,1653,303);
  `device_slave_connections_TB_CONFIG_4(2,1654,304);
  `device_slave_connections_TB_CONFIG_4(2,1655,305);
  `device_slave_connections_TB_CONFIG_4(2,1656,306);
  `device_slave_connections_TB_CONFIG_4(2,1657,307);
  `device_slave_connections_TB_CONFIG_4(2,1658,308);
  `device_slave_connections_TB_CONFIG_4(2,1659,309);
  `device_slave_connections_TB_CONFIG_4(2,1660,310);
  `device_slave_connections_TB_CONFIG_4(2,1661,311);
  `device_slave_connections_TB_CONFIG_4(2,1662,312);
  `device_slave_connections_TB_CONFIG_4(2,1663,313);
  `device_slave_connections_TB_CONFIG_4(2,1664,314);
  `device_slave_connections_TB_CONFIG_4(2,1665,315);
  `device_slave_connections_TB_CONFIG_4(2,1666,316);
  `device_slave_connections_TB_CONFIG_4(2,1667,317);
  `device_slave_connections_TB_CONFIG_4(2,1668,318);
  `device_slave_connections_TB_CONFIG_4(2,1669,319);
  `device_slave_connections_TB_CONFIG_4(2,1670,320);
  `device_slave_connections_TB_CONFIG_4(2,1671,321);
  `device_slave_connections_TB_CONFIG_4(2,1672,322);
  `device_slave_connections_TB_CONFIG_4(2,1673,323);
  `device_slave_connections_TB_CONFIG_4(2,1674,324);
  `device_slave_connections_TB_CONFIG_4(2,1675,325);
  `device_slave_connections_TB_CONFIG_4(2,1676,326);
  `device_slave_connections_TB_CONFIG_4(2,1677,327);
  `device_slave_connections_TB_CONFIG_4(2,1678,328);
  `device_slave_connections_TB_CONFIG_4(2,1679,329);
  `device_slave_connections_TB_CONFIG_4(2,1680,330);
  `device_slave_connections_TB_CONFIG_4(2,1681,331);
  `device_slave_connections_TB_CONFIG_4(2,1682,332);
  `device_slave_connections_TB_CONFIG_4(2,1683,333);
  `device_slave_connections_TB_CONFIG_4(2,1684,334);
  `device_slave_connections_TB_CONFIG_4(2,1685,335);
  `device_slave_connections_TB_CONFIG_4(2,1686,336);
  `device_slave_connections_TB_CONFIG_4(2,1687,337);
  `device_slave_connections_TB_CONFIG_4(2,1688,338);
  `device_slave_connections_TB_CONFIG_4(2,1689,339);
  `device_slave_connections_TB_CONFIG_4(2,1690,340);
  `device_slave_connections_TB_CONFIG_4(2,1691,341);
  `device_slave_connections_TB_CONFIG_4(2,1692,342);
  `device_slave_connections_TB_CONFIG_4(2,1693,343);
  `device_slave_connections_TB_CONFIG_4(2,1694,344);
  `device_slave_connections_TB_CONFIG_4(2,1695,345);
  `device_slave_connections_TB_CONFIG_4(2,1696,346);
  `device_slave_connections_TB_CONFIG_4(2,1697,347);
  `device_slave_connections_TB_CONFIG_4(2,1698,348);
  `device_slave_connections_TB_CONFIG_4(2,1699,349);
  `device_slave_connections_TB_CONFIG_4(2,1700,350);
  `device_slave_connections_TB_CONFIG_4(2,1701,351);
  `device_slave_connections_TB_CONFIG_4(2,1702,352);
  `device_slave_connections_TB_CONFIG_4(2,1703,353);
  `device_slave_connections_TB_CONFIG_4(2,1704,354);
  `device_slave_connections_TB_CONFIG_4(2,1705,355);
  `device_slave_connections_TB_CONFIG_4(2,1706,356);
  `device_slave_connections_TB_CONFIG_4(2,1707,357);
  `device_slave_connections_TB_CONFIG_4(2,1708,358);
  `device_slave_connections_TB_CONFIG_4(2,1709,359);
  `device_slave_connections_TB_CONFIG_4(2,1710,360);
  `device_slave_connections_TB_CONFIG_4(2,1711,361);
  `device_slave_connections_TB_CONFIG_4(2,1712,362);
  `device_slave_connections_TB_CONFIG_4(2,1713,363);
  `device_slave_connections_TB_CONFIG_4(2,1714,364);
  `device_slave_connections_TB_CONFIG_4(2,1715,365);
  `device_slave_connections_TB_CONFIG_4(2,1716,366);
  `device_slave_connections_TB_CONFIG_4(2,1717,367);
  `device_slave_connections_TB_CONFIG_4(2,1718,368);
  `device_slave_connections_TB_CONFIG_4(2,1719,369);
  `device_slave_connections_TB_CONFIG_4(2,1720,370);
  `device_slave_connections_TB_CONFIG_4(2,1721,371);
  `device_slave_connections_TB_CONFIG_4(2,1722,372);
  `device_slave_connections_TB_CONFIG_4(2,1723,373);
  `device_slave_connections_TB_CONFIG_4(2,1724,374);
  `device_slave_connections_TB_CONFIG_4(2,1725,375);
  `device_slave_connections_TB_CONFIG_4(2,1726,376);
  `device_slave_connections_TB_CONFIG_4(2,1727,377);
  `device_slave_connections_TB_CONFIG_4(2,1728,378);
  `device_slave_connections_TB_CONFIG_4(2,1729,379);
  `device_slave_connections_TB_CONFIG_4(2,1730,380);
  `device_slave_connections_TB_CONFIG_4(2,1731,381);
  `device_slave_connections_TB_CONFIG_4(2,1732,382);
  `device_slave_connections_TB_CONFIG_4(2,1733,383);
  `device_slave_connections_TB_CONFIG_4(2,1734,384);
  `device_slave_connections_TB_CONFIG_4(2,1735,385);
  `device_slave_connections_TB_CONFIG_4(2,1736,386);
  `device_slave_connections_TB_CONFIG_4(2,1737,387);
  `device_slave_connections_TB_CONFIG_4(2,1738,388);
  `device_slave_connections_TB_CONFIG_4(2,1739,389);
  `device_slave_connections_TB_CONFIG_4(2,1740,390);
  `device_slave_connections_TB_CONFIG_4(2,1741,391);
  `device_slave_connections_TB_CONFIG_4(2,1742,392);
  `device_slave_connections_TB_CONFIG_4(2,1743,393);
  `device_slave_connections_TB_CONFIG_4(2,1744,394);
  `device_slave_connections_TB_CONFIG_4(2,1745,395);
  `device_slave_connections_TB_CONFIG_4(2,1746,396);
  `device_slave_connections_TB_CONFIG_4(2,1747,397);
  `device_slave_connections_TB_CONFIG_4(2,1748,398);
  `device_slave_connections_TB_CONFIG_4(2,1749,399);
  `device_slave_connections_TB_CONFIG_4(2,1750,400);
  `device_slave_connections_TB_CONFIG_4(2,1751,401);
  `device_slave_connections_TB_CONFIG_4(2,1752,402);
  `device_slave_connections_TB_CONFIG_4(2,1753,403);
  `device_slave_connections_TB_CONFIG_4(2,1754,404);
  `device_slave_connections_TB_CONFIG_4(2,1755,405);
  `device_slave_connections_TB_CONFIG_4(2,1756,406);
  `device_slave_connections_TB_CONFIG_4(2,1757,407);
  `device_slave_connections_TB_CONFIG_4(2,1758,408);
  `device_slave_connections_TB_CONFIG_4(2,1759,409);
  `device_slave_connections_TB_CONFIG_4(2,1760,410);
  `device_slave_connections_TB_CONFIG_4(2,1761,411);
  `device_slave_connections_TB_CONFIG_4(2,1762,412);
  `device_slave_connections_TB_CONFIG_4(2,1763,413);
  `device_slave_connections_TB_CONFIG_4(2,1764,414);
  `device_slave_connections_TB_CONFIG_4(2,1765,415);
  `device_slave_connections_TB_CONFIG_4(2,1766,416);
  `device_slave_connections_TB_CONFIG_4(2,1767,417);
  `device_slave_connections_TB_CONFIG_4(2,1768,418);
  `device_slave_connections_TB_CONFIG_4(2,1769,419);
  `device_slave_connections_TB_CONFIG_4(2,1770,420);
  `device_slave_connections_TB_CONFIG_4(2,1771,421);
  `device_slave_connections_TB_CONFIG_4(2,1772,422);
  `device_slave_connections_TB_CONFIG_4(2,1773,423);
  `device_slave_connections_TB_CONFIG_4(2,1774,424);
  `device_slave_connections_TB_CONFIG_4(2,1775,425);
  `device_slave_connections_TB_CONFIG_4(2,1776,426);
  `device_slave_connections_TB_CONFIG_4(2,1777,427);
  `device_slave_connections_TB_CONFIG_4(2,1778,428);
  `device_slave_connections_TB_CONFIG_4(2,1779,429);
  `device_slave_connections_TB_CONFIG_4(2,1780,430);
  `device_slave_connections_TB_CONFIG_4(2,1781,431);
  `device_slave_connections_TB_CONFIG_4(2,1782,432);
  `device_slave_connections_TB_CONFIG_4(2,1783,433);
  `device_slave_connections_TB_CONFIG_4(2,1784,434);
  `device_slave_connections_TB_CONFIG_4(2,1785,435);
  `device_slave_connections_TB_CONFIG_4(2,1786,436);
  `device_slave_connections_TB_CONFIG_4(2,1787,437);
  `device_slave_connections_TB_CONFIG_4(2,1788,438);
  `device_slave_connections_TB_CONFIG_4(2,1789,439);
  `device_slave_connections_TB_CONFIG_4(2,1790,440);
  `device_slave_connections_TB_CONFIG_4(2,1791,441);
  `device_slave_connections_TB_CONFIG_4(2,1792,442);
  `device_slave_connections_TB_CONFIG_4(2,1793,443);
  `device_slave_connections_TB_CONFIG_4(2,1794,444);
  `device_slave_connections_TB_CONFIG_4(2,1795,445);
  `device_slave_connections_TB_CONFIG_4(2,1796,446);
  `device_slave_connections_TB_CONFIG_4(2,1797,447);
  `device_slave_connections_TB_CONFIG_4(2,1798,448);
  `device_slave_connections_TB_CONFIG_4(2,1799,449);
	`device_slave_connections_TB_CONFIG_4(3,1800,0);
  `device_slave_connections_TB_CONFIG_4(3,1801,1);
  `device_slave_connections_TB_CONFIG_4(3,1802,2);
  `device_slave_connections_TB_CONFIG_4(3,1803,3);
  `device_slave_connections_TB_CONFIG_4(3,1804,4);
  `device_slave_connections_TB_CONFIG_4(3,1805,5);
  `device_slave_connections_TB_CONFIG_4(3,1806,6);
  `device_slave_connections_TB_CONFIG_4(3,1807,7);
  `device_slave_connections_TB_CONFIG_4(3,1808,8);
  `device_slave_connections_TB_CONFIG_4(3,1809,9);
  `device_slave_connections_TB_CONFIG_4(3,1810,10);
  `device_slave_connections_TB_CONFIG_4(3,1811,11);
  `device_slave_connections_TB_CONFIG_4(3,1812,12);
  `device_slave_connections_TB_CONFIG_4(3,1813,13);
  `device_slave_connections_TB_CONFIG_4(3,1814,14);
  `device_slave_connections_TB_CONFIG_4(3,1815,15);
  `device_slave_connections_TB_CONFIG_4(3,1816,16);
  `device_slave_connections_TB_CONFIG_4(3,1817,17);
  `device_slave_connections_TB_CONFIG_4(3,1818,18);
  `device_slave_connections_TB_CONFIG_4(3,1819,19);
  `device_slave_connections_TB_CONFIG_4(3,1820,20);
  `device_slave_connections_TB_CONFIG_4(3,1821,21);
  `device_slave_connections_TB_CONFIG_4(3,1822,22);
  `device_slave_connections_TB_CONFIG_4(3,1823,23);
  `device_slave_connections_TB_CONFIG_4(3,1824,24);
  `device_slave_connections_TB_CONFIG_4(3,1825,25);
  `device_slave_connections_TB_CONFIG_4(3,1826,26);
  `device_slave_connections_TB_CONFIG_4(3,1827,27);
  `device_slave_connections_TB_CONFIG_4(3,1828,28);
  `device_slave_connections_TB_CONFIG_4(3,1829,29);
  `device_slave_connections_TB_CONFIG_4(3,1830,30);
  `device_slave_connections_TB_CONFIG_4(3,1831,31);
  `device_slave_connections_TB_CONFIG_4(3,1832,32);
  `device_slave_connections_TB_CONFIG_4(3,1833,33);
  `device_slave_connections_TB_CONFIG_4(3,1834,34);
  `device_slave_connections_TB_CONFIG_4(3,1835,35);
  `device_slave_connections_TB_CONFIG_4(3,1836,36);
  `device_slave_connections_TB_CONFIG_4(3,1837,37);
  `device_slave_connections_TB_CONFIG_4(3,1838,38);
  `device_slave_connections_TB_CONFIG_4(3,1839,39);
  `device_slave_connections_TB_CONFIG_4(3,1840,40);
  `device_slave_connections_TB_CONFIG_4(3,1841,41);
  `device_slave_connections_TB_CONFIG_4(3,1842,42);
  `device_slave_connections_TB_CONFIG_4(3,1843,43);
  `device_slave_connections_TB_CONFIG_4(3,1844,44);
  `device_slave_connections_TB_CONFIG_4(3,1845,45);
  `device_slave_connections_TB_CONFIG_4(3,1846,46);
  `device_slave_connections_TB_CONFIG_4(3,1847,47);
  `device_slave_connections_TB_CONFIG_4(3,1848,48);
  `device_slave_connections_TB_CONFIG_4(3,1849,49);
  `device_slave_connections_TB_CONFIG_4(3,1850,50);
  `device_slave_connections_TB_CONFIG_4(3,1851,51);
  `device_slave_connections_TB_CONFIG_4(3,1852,52);
  `device_slave_connections_TB_CONFIG_4(3,1853,53);
  `device_slave_connections_TB_CONFIG_4(3,1854,54);
  `device_slave_connections_TB_CONFIG_4(3,1855,55);
  `device_slave_connections_TB_CONFIG_4(3,1856,56);
  `device_slave_connections_TB_CONFIG_4(3,1857,57);
  `device_slave_connections_TB_CONFIG_4(3,1858,58);
  `device_slave_connections_TB_CONFIG_4(3,1859,59);
  `device_slave_connections_TB_CONFIG_4(3,1860,60);
  `device_slave_connections_TB_CONFIG_4(3,1861,61);
  `device_slave_connections_TB_CONFIG_4(3,1862,62);
  `device_slave_connections_TB_CONFIG_4(3,1863,63);
  `device_slave_connections_TB_CONFIG_4(3,1864,64);
  `device_slave_connections_TB_CONFIG_4(3,1865,65);
  `device_slave_connections_TB_CONFIG_4(3,1866,66);
  `device_slave_connections_TB_CONFIG_4(3,1867,67);
  `device_slave_connections_TB_CONFIG_4(3,1868,68);
  `device_slave_connections_TB_CONFIG_4(3,1869,69);
  `device_slave_connections_TB_CONFIG_4(3,1870,70);
  `device_slave_connections_TB_CONFIG_4(3,1871,71);
  `device_slave_connections_TB_CONFIG_4(3,1872,72);
  `device_slave_connections_TB_CONFIG_4(3,1873,73);
  `device_slave_connections_TB_CONFIG_4(3,1874,74);
  `device_slave_connections_TB_CONFIG_4(3,1875,75);
  `device_slave_connections_TB_CONFIG_4(3,1876,76);
  `device_slave_connections_TB_CONFIG_4(3,1877,77);
  `device_slave_connections_TB_CONFIG_4(3,1878,78);
  `device_slave_connections_TB_CONFIG_4(3,1879,79);
  `device_slave_connections_TB_CONFIG_4(3,1880,80);
  `device_slave_connections_TB_CONFIG_4(3,1881,81);
  `device_slave_connections_TB_CONFIG_4(3,1882,82);
  `device_slave_connections_TB_CONFIG_4(3,1883,83);
  `device_slave_connections_TB_CONFIG_4(3,1884,84);
  `device_slave_connections_TB_CONFIG_4(3,1885,85);
  `device_slave_connections_TB_CONFIG_4(3,1886,86);
  `device_slave_connections_TB_CONFIG_4(3,1887,87);
  `device_slave_connections_TB_CONFIG_4(3,1888,88);
  `device_slave_connections_TB_CONFIG_4(3,1889,89);
  `device_slave_connections_TB_CONFIG_4(3,1890,90);
  `device_slave_connections_TB_CONFIG_4(3,1891,91);
  `device_slave_connections_TB_CONFIG_4(3,1892,92);
  `device_slave_connections_TB_CONFIG_4(3,1893,93);
  `device_slave_connections_TB_CONFIG_4(3,1894,94);
  `device_slave_connections_TB_CONFIG_4(3,1895,95);
  `device_slave_connections_TB_CONFIG_4(3,1896,96);
  `device_slave_connections_TB_CONFIG_4(3,1897,97);
  `device_slave_connections_TB_CONFIG_4(3,1898,98);
  `device_slave_connections_TB_CONFIG_4(3,1899,99);
  `device_slave_connections_TB_CONFIG_4(3,1900,100);
  `device_slave_connections_TB_CONFIG_4(3,1901,101);
  `device_slave_connections_TB_CONFIG_4(3,1902,102);
  `device_slave_connections_TB_CONFIG_4(3,1903,103);
  `device_slave_connections_TB_CONFIG_4(3,1904,104);
  `device_slave_connections_TB_CONFIG_4(3,1905,105);
  `device_slave_connections_TB_CONFIG_4(3,1906,106);
  `device_slave_connections_TB_CONFIG_4(3,1907,107);
  `device_slave_connections_TB_CONFIG_4(3,1908,108);
  `device_slave_connections_TB_CONFIG_4(3,1909,109);
  `device_slave_connections_TB_CONFIG_4(3,1910,110);
  `device_slave_connections_TB_CONFIG_4(3,1911,111);
  `device_slave_connections_TB_CONFIG_4(3,1912,112);
  `device_slave_connections_TB_CONFIG_4(3,1913,113);
  `device_slave_connections_TB_CONFIG_4(3,1914,114);
  `device_slave_connections_TB_CONFIG_4(3,1915,115);
  `device_slave_connections_TB_CONFIG_4(3,1916,116);
  `device_slave_connections_TB_CONFIG_4(3,1917,117);
  `device_slave_connections_TB_CONFIG_4(3,1918,118);
  `device_slave_connections_TB_CONFIG_4(3,1919,119);
  `device_slave_connections_TB_CONFIG_4(3,1920,120);
  `device_slave_connections_TB_CONFIG_4(3,1921,121);
  `device_slave_connections_TB_CONFIG_4(3,1922,122);
  `device_slave_connections_TB_CONFIG_4(3,1923,123);
  `device_slave_connections_TB_CONFIG_4(3,1924,124);
  `device_slave_connections_TB_CONFIG_4(3,1925,125);
  `device_slave_connections_TB_CONFIG_4(3,1926,126);
  `device_slave_connections_TB_CONFIG_4(3,1927,127);
  `device_slave_connections_TB_CONFIG_4(3,1928,128);
  `device_slave_connections_TB_CONFIG_4(3,1929,129);
  `device_slave_connections_TB_CONFIG_4(3,1930,130);
  `device_slave_connections_TB_CONFIG_4(3,1931,131);
  `device_slave_connections_TB_CONFIG_4(3,1932,132);
  `device_slave_connections_TB_CONFIG_4(3,1933,133);
  `device_slave_connections_TB_CONFIG_4(3,1934,134);
  `device_slave_connections_TB_CONFIG_4(3,1935,135);
  `device_slave_connections_TB_CONFIG_4(3,1936,136);
  `device_slave_connections_TB_CONFIG_4(3,1937,137);
  `device_slave_connections_TB_CONFIG_4(3,1938,138);
  `device_slave_connections_TB_CONFIG_4(3,1939,139);
  `device_slave_connections_TB_CONFIG_4(3,1940,140);
  `device_slave_connections_TB_CONFIG_4(3,1941,141);
  `device_slave_connections_TB_CONFIG_4(3,1942,142);
  `device_slave_connections_TB_CONFIG_4(3,1943,143);
  `device_slave_connections_TB_CONFIG_4(3,1944,144);
  `device_slave_connections_TB_CONFIG_4(3,1945,145);
  `device_slave_connections_TB_CONFIG_4(3,1946,146);
  `device_slave_connections_TB_CONFIG_4(3,1947,147);
  `device_slave_connections_TB_CONFIG_4(3,1948,148);
  `device_slave_connections_TB_CONFIG_4(3,1949,149);
  `device_slave_connections_TB_CONFIG_4(3,1950,150);
  `device_slave_connections_TB_CONFIG_4(3,1951,151);
  `device_slave_connections_TB_CONFIG_4(3,1952,152);
  `device_slave_connections_TB_CONFIG_4(3,1953,153);
  `device_slave_connections_TB_CONFIG_4(3,1954,154);
  `device_slave_connections_TB_CONFIG_4(3,1955,155);
  `device_slave_connections_TB_CONFIG_4(3,1956,156);
  `device_slave_connections_TB_CONFIG_4(3,1957,157);
  `device_slave_connections_TB_CONFIG_4(3,1958,158);
  `device_slave_connections_TB_CONFIG_4(3,1959,159);
  `device_slave_connections_TB_CONFIG_4(3,1960,160);
  `device_slave_connections_TB_CONFIG_4(3,1961,161);
  `device_slave_connections_TB_CONFIG_4(3,1962,162);
  `device_slave_connections_TB_CONFIG_4(3,1963,163);
  `device_slave_connections_TB_CONFIG_4(3,1964,164);
  `device_slave_connections_TB_CONFIG_4(3,1965,165);
  `device_slave_connections_TB_CONFIG_4(3,1966,166);
  `device_slave_connections_TB_CONFIG_4(3,1967,167);
  `device_slave_connections_TB_CONFIG_4(3,1968,168);
  `device_slave_connections_TB_CONFIG_4(3,1969,169);
  `device_slave_connections_TB_CONFIG_4(3,1970,170);
  `device_slave_connections_TB_CONFIG_4(3,1971,171);
  `device_slave_connections_TB_CONFIG_4(3,1972,172);
  `device_slave_connections_TB_CONFIG_4(3,1973,173);
  `device_slave_connections_TB_CONFIG_4(3,1974,174);
  `device_slave_connections_TB_CONFIG_4(3,1975,175);
  `device_slave_connections_TB_CONFIG_4(3,1976,176);
  `device_slave_connections_TB_CONFIG_4(3,1977,177);
  `device_slave_connections_TB_CONFIG_4(3,1978,178);
  `device_slave_connections_TB_CONFIG_4(3,1979,179);
  `device_slave_connections_TB_CONFIG_4(3,1980,180);
  `device_slave_connections_TB_CONFIG_4(3,1981,181);
  `device_slave_connections_TB_CONFIG_4(3,1982,182);
  `device_slave_connections_TB_CONFIG_4(3,1983,183);
  `device_slave_connections_TB_CONFIG_4(3,1984,184);
  `device_slave_connections_TB_CONFIG_4(3,1985,185);
  `device_slave_connections_TB_CONFIG_4(3,1986,186);
  `device_slave_connections_TB_CONFIG_4(3,1987,187);
  `device_slave_connections_TB_CONFIG_4(3,1988,188);
  `device_slave_connections_TB_CONFIG_4(3,1989,189);
  `device_slave_connections_TB_CONFIG_4(3,1990,190);
  `device_slave_connections_TB_CONFIG_4(3,1991,191);
  `device_slave_connections_TB_CONFIG_4(3,1992,192);
  `device_slave_connections_TB_CONFIG_4(3,1993,193);
  `device_slave_connections_TB_CONFIG_4(3,1994,194);
  `device_slave_connections_TB_CONFIG_4(3,1995,195);
  `device_slave_connections_TB_CONFIG_4(3,1996,196);
  `device_slave_connections_TB_CONFIG_4(3,1997,197);
  `device_slave_connections_TB_CONFIG_4(3,1998,198);
  `device_slave_connections_TB_CONFIG_4(3,1999,199);
  `device_slave_connections_TB_CONFIG_4(3,2000,200);
  `device_slave_connections_TB_CONFIG_4(3,2001,201);
  `device_slave_connections_TB_CONFIG_4(3,2002,202);
  `device_slave_connections_TB_CONFIG_4(3,2003,203);
  `device_slave_connections_TB_CONFIG_4(3,2004,204);
  `device_slave_connections_TB_CONFIG_4(3,2005,205);
  `device_slave_connections_TB_CONFIG_4(3,2006,206);
  `device_slave_connections_TB_CONFIG_4(3,2007,207);
  `device_slave_connections_TB_CONFIG_4(3,2008,208);
  `device_slave_connections_TB_CONFIG_4(3,2009,209);
  `device_slave_connections_TB_CONFIG_4(3,2010,210);
  `device_slave_connections_TB_CONFIG_4(3,2011,211);
  `device_slave_connections_TB_CONFIG_4(3,2012,212);
  `device_slave_connections_TB_CONFIG_4(3,2013,213);
  `device_slave_connections_TB_CONFIG_4(3,2014,214);
  `device_slave_connections_TB_CONFIG_4(3,2015,215);
  `device_slave_connections_TB_CONFIG_4(3,2016,216);
  `device_slave_connections_TB_CONFIG_4(3,2017,217);
  `device_slave_connections_TB_CONFIG_4(3,2018,218);
  `device_slave_connections_TB_CONFIG_4(3,2019,219);
  `device_slave_connections_TB_CONFIG_4(3,2020,220);
  `device_slave_connections_TB_CONFIG_4(3,2021,221);
  `device_slave_connections_TB_CONFIG_4(3,2022,222);
  `device_slave_connections_TB_CONFIG_4(3,2023,223);
  `device_slave_connections_TB_CONFIG_4(3,2024,224);
  `device_slave_connections_TB_CONFIG_4(3,2025,225);
  `device_slave_connections_TB_CONFIG_4(3,2026,226);
  `device_slave_connections_TB_CONFIG_4(3,2027,227);
  `device_slave_connections_TB_CONFIG_4(3,2028,228);
  `device_slave_connections_TB_CONFIG_4(3,2029,229);
  `device_slave_connections_TB_CONFIG_4(3,2030,230);
  `device_slave_connections_TB_CONFIG_4(3,2031,231);
  `device_slave_connections_TB_CONFIG_4(3,2032,232);
  `device_slave_connections_TB_CONFIG_4(3,2033,233);
  `device_slave_connections_TB_CONFIG_4(3,2034,234);
  `device_slave_connections_TB_CONFIG_4(3,2035,235);
  `device_slave_connections_TB_CONFIG_4(3,2036,236);
  `device_slave_connections_TB_CONFIG_4(3,2037,237);
  `device_slave_connections_TB_CONFIG_4(3,2038,238);
  `device_slave_connections_TB_CONFIG_4(3,2039,239);
  `device_slave_connections_TB_CONFIG_4(3,2040,240);
  `device_slave_connections_TB_CONFIG_4(3,2041,241);
  `device_slave_connections_TB_CONFIG_4(3,2042,242);
  `device_slave_connections_TB_CONFIG_4(3,2043,243);
  `device_slave_connections_TB_CONFIG_4(3,2044,244);
  `device_slave_connections_TB_CONFIG_4(3,2045,245);
  `device_slave_connections_TB_CONFIG_4(3,2046,246);
  `device_slave_connections_TB_CONFIG_4(3,2047,247);
  /*`device_slave_connections_TB_CONFIG_4(3,2048,248);
  `device_slave_connections_TB_CONFIG_4(3,2049,249);
  `device_slave_connections_TB_CONFIG_4(3,2050,250);
  `device_slave_connections_TB_CONFIG_4(3,2051,251);
  `device_slave_connections_TB_CONFIG_4(3,2052,252);
  `device_slave_connections_TB_CONFIG_4(3,2053,253);
  `device_slave_connections_TB_CONFIG_4(3,2054,254);
  `device_slave_connections_TB_CONFIG_4(3,2055,255);
  `device_slave_connections_TB_CONFIG_4(3,2056,256);
  `device_slave_connections_TB_CONFIG_4(3,2057,257);
  `device_slave_connections_TB_CONFIG_4(3,2058,258);
  `device_slave_connections_TB_CONFIG_4(3,2059,259);
  `device_slave_connections_TB_CONFIG_4(3,2060,260);
  `device_slave_connections_TB_CONFIG_4(3,2061,261);
  `device_slave_connections_TB_CONFIG_4(3,2062,262);
  `device_slave_connections_TB_CONFIG_4(3,2063,263);
  `device_slave_connections_TB_CONFIG_4(3,2064,264);
  `device_slave_connections_TB_CONFIG_4(3,2065,265);
  `device_slave_connections_TB_CONFIG_4(3,2066,266);
  `device_slave_connections_TB_CONFIG_4(3,2067,267);
  `device_slave_connections_TB_CONFIG_4(3,2068,268);
  `device_slave_connections_TB_CONFIG_4(3,2069,269);
  `device_slave_connections_TB_CONFIG_4(3,2070,270);
  `device_slave_connections_TB_CONFIG_4(3,2071,271);
  `device_slave_connections_TB_CONFIG_4(3,2072,272);
  `device_slave_connections_TB_CONFIG_4(3,2073,273);
  `device_slave_connections_TB_CONFIG_4(3,2074,274);
  `device_slave_connections_TB_CONFIG_4(3,2075,275);
  `device_slave_connections_TB_CONFIG_4(3,2076,276);
  `device_slave_connections_TB_CONFIG_4(3,2077,277);
  `device_slave_connections_TB_CONFIG_4(3,2078,278);
  `device_slave_connections_TB_CONFIG_4(3,2079,279);
  `device_slave_connections_TB_CONFIG_4(3,2080,280);
  `device_slave_connections_TB_CONFIG_4(3,2081,281);
  `device_slave_connections_TB_CONFIG_4(3,2082,282);
  `device_slave_connections_TB_CONFIG_4(3,2083,283);
  `device_slave_connections_TB_CONFIG_4(3,2084,284);
  `device_slave_connections_TB_CONFIG_4(3,2085,285);
  `device_slave_connections_TB_CONFIG_4(3,2086,286);
  `device_slave_connections_TB_CONFIG_4(3,2087,287);
  `device_slave_connections_TB_CONFIG_4(3,2088,288);
  `device_slave_connections_TB_CONFIG_4(3,2089,289);
  `device_slave_connections_TB_CONFIG_4(3,2090,290);
  `device_slave_connections_TB_CONFIG_4(3,2091,291);
  `device_slave_connections_TB_CONFIG_4(3,2092,292);
  `device_slave_connections_TB_CONFIG_4(3,2093,293);
  `device_slave_connections_TB_CONFIG_4(3,2094,294);
  `device_slave_connections_TB_CONFIG_4(3,2095,295);
  `device_slave_connections_TB_CONFIG_4(3,2096,296);
  `device_slave_connections_TB_CONFIG_4(3,2097,297);
  `device_slave_connections_TB_CONFIG_4(3,2098,298);
  `device_slave_connections_TB_CONFIG_4(3,2099,299);
  `device_slave_connections_TB_CONFIG_4(3,2100,300);
  `device_slave_connections_TB_CONFIG_4(3,2101,301);
  `device_slave_connections_TB_CONFIG_4(3,2102,302);
  `device_slave_connections_TB_CONFIG_4(3,2103,303);
  `device_slave_connections_TB_CONFIG_4(3,2104,304);
  `device_slave_connections_TB_CONFIG_4(3,2105,305);
  `device_slave_connections_TB_CONFIG_4(3,2106,306);
  `device_slave_connections_TB_CONFIG_4(3,2107,307);
  `device_slave_connections_TB_CONFIG_4(3,2108,308);
  `device_slave_connections_TB_CONFIG_4(3,2109,309);
  `device_slave_connections_TB_CONFIG_4(3,2110,310);
  `device_slave_connections_TB_CONFIG_4(3,2111,311);
  `device_slave_connections_TB_CONFIG_4(3,2112,312);
  `device_slave_connections_TB_CONFIG_4(3,2113,313);
  `device_slave_connections_TB_CONFIG_4(3,2114,314);
  `device_slave_connections_TB_CONFIG_4(3,2115,315);
  `device_slave_connections_TB_CONFIG_4(3,2116,316);
  `device_slave_connections_TB_CONFIG_4(3,2117,317);
  `device_slave_connections_TB_CONFIG_4(3,2118,318);
  `device_slave_connections_TB_CONFIG_4(3,2119,319);
  `device_slave_connections_TB_CONFIG_4(3,2120,320);
  `device_slave_connections_TB_CONFIG_4(3,2121,321);
  `device_slave_connections_TB_CONFIG_4(3,2122,322);
  `device_slave_connections_TB_CONFIG_4(3,2123,323);
  `device_slave_connections_TB_CONFIG_4(3,2124,324);
  `device_slave_connections_TB_CONFIG_4(3,2125,325);
  `device_slave_connections_TB_CONFIG_4(3,2126,326);
  `device_slave_connections_TB_CONFIG_4(3,2127,327);
  `device_slave_connections_TB_CONFIG_4(3,2128,328);
  `device_slave_connections_TB_CONFIG_4(3,2129,329);
  `device_slave_connections_TB_CONFIG_4(3,2130,330);
  `device_slave_connections_TB_CONFIG_4(3,2131,331);
  `device_slave_connections_TB_CONFIG_4(3,2132,332);
  `device_slave_connections_TB_CONFIG_4(3,2133,333);
  `device_slave_connections_TB_CONFIG_4(3,2134,334);
  `device_slave_connections_TB_CONFIG_4(3,2135,335);
  `device_slave_connections_TB_CONFIG_4(3,2136,336);
  `device_slave_connections_TB_CONFIG_4(3,2137,337);
  `device_slave_connections_TB_CONFIG_4(3,2138,338);
  `device_slave_connections_TB_CONFIG_4(3,2139,339);
  `device_slave_connections_TB_CONFIG_4(3,2140,340);
  `device_slave_connections_TB_CONFIG_4(3,2141,341);
  `device_slave_connections_TB_CONFIG_4(3,2142,342);
  `device_slave_connections_TB_CONFIG_4(3,2143,343);
  `device_slave_connections_TB_CONFIG_4(3,2144,344);
  `device_slave_connections_TB_CONFIG_4(3,2145,345);
  `device_slave_connections_TB_CONFIG_4(3,2146,346);
  `device_slave_connections_TB_CONFIG_4(3,2147,347);
  `device_slave_connections_TB_CONFIG_4(3,2148,348);
  `device_slave_connections_TB_CONFIG_4(3,2149,349);
  `device_slave_connections_TB_CONFIG_4(3,2150,350);
  `device_slave_connections_TB_CONFIG_4(3,2151,351);
  `device_slave_connections_TB_CONFIG_4(3,2152,352);
  `device_slave_connections_TB_CONFIG_4(3,2153,353);
  `device_slave_connections_TB_CONFIG_4(3,2154,354);
  `device_slave_connections_TB_CONFIG_4(3,2155,355);
  `device_slave_connections_TB_CONFIG_4(3,2156,356);
  `device_slave_connections_TB_CONFIG_4(3,2157,357);
  `device_slave_connections_TB_CONFIG_4(3,2158,358);
  `device_slave_connections_TB_CONFIG_4(3,2159,359);
  `device_slave_connections_TB_CONFIG_4(3,2160,360);
  `device_slave_connections_TB_CONFIG_4(3,2161,361);
  `device_slave_connections_TB_CONFIG_4(3,2162,362);
  `device_slave_connections_TB_CONFIG_4(3,2163,363);
  `device_slave_connections_TB_CONFIG_4(3,2164,364);
  `device_slave_connections_TB_CONFIG_4(3,2165,365);
  `device_slave_connections_TB_CONFIG_4(3,2166,366);
  `device_slave_connections_TB_CONFIG_4(3,2167,367);
  `device_slave_connections_TB_CONFIG_4(3,2168,368);
  `device_slave_connections_TB_CONFIG_4(3,2169,369);
  `device_slave_connections_TB_CONFIG_4(3,2170,370);
  `device_slave_connections_TB_CONFIG_4(3,2171,371);
  `device_slave_connections_TB_CONFIG_4(3,2172,372);
  `device_slave_connections_TB_CONFIG_4(3,2173,373);
  `device_slave_connections_TB_CONFIG_4(3,2174,374);
  `device_slave_connections_TB_CONFIG_4(3,2175,375);
  `device_slave_connections_TB_CONFIG_4(3,2176,376);
  `device_slave_connections_TB_CONFIG_4(3,2177,377);
  `device_slave_connections_TB_CONFIG_4(3,2178,378);
  `device_slave_connections_TB_CONFIG_4(3,2179,379);
  `device_slave_connections_TB_CONFIG_4(3,2180,380);
  `device_slave_connections_TB_CONFIG_4(3,2181,381);
  `device_slave_connections_TB_CONFIG_4(3,2182,382);
  `device_slave_connections_TB_CONFIG_4(3,2183,383);
  `device_slave_connections_TB_CONFIG_4(3,2184,384);
  `device_slave_connections_TB_CONFIG_4(3,2185,385);
  `device_slave_connections_TB_CONFIG_4(3,2186,386);
  `device_slave_connections_TB_CONFIG_4(3,2187,387);
  `device_slave_connections_TB_CONFIG_4(3,2188,388);
  `device_slave_connections_TB_CONFIG_4(3,2189,389);
  `device_slave_connections_TB_CONFIG_4(3,2190,390);
  `device_slave_connections_TB_CONFIG_4(3,2191,391);
  `device_slave_connections_TB_CONFIG_4(3,2192,392);
  `device_slave_connections_TB_CONFIG_4(3,2193,393);
  `device_slave_connections_TB_CONFIG_4(3,2194,394);
  `device_slave_connections_TB_CONFIG_4(3,2195,395);
  `device_slave_connections_TB_CONFIG_4(3,2196,396);
  `device_slave_connections_TB_CONFIG_4(3,2197,397);
  `device_slave_connections_TB_CONFIG_4(3,2198,398);
  `device_slave_connections_TB_CONFIG_4(3,2199,399);
  `device_slave_connections_TB_CONFIG_4(3,2200,400);
  `device_slave_connections_TB_CONFIG_4(3,2201,401);
  `device_slave_connections_TB_CONFIG_4(3,2202,402);
  `device_slave_connections_TB_CONFIG_4(3,2203,403);
  `device_slave_connections_TB_CONFIG_4(3,2204,404);
  `device_slave_connections_TB_CONFIG_4(3,2205,405);
  `device_slave_connections_TB_CONFIG_4(3,2206,406);
  `device_slave_connections_TB_CONFIG_4(3,2207,407);
  `device_slave_connections_TB_CONFIG_4(3,2208,408);
  `device_slave_connections_TB_CONFIG_4(3,2209,409);
  `device_slave_connections_TB_CONFIG_4(3,2210,410);
  `device_slave_connections_TB_CONFIG_4(3,2211,411);
  `device_slave_connections_TB_CONFIG_4(3,2212,412);
  `device_slave_connections_TB_CONFIG_4(3,2213,413);
  `device_slave_connections_TB_CONFIG_4(3,2214,414);
  `device_slave_connections_TB_CONFIG_4(3,2215,415);
  `device_slave_connections_TB_CONFIG_4(3,2216,416);
  `device_slave_connections_TB_CONFIG_4(3,2217,417);
  `device_slave_connections_TB_CONFIG_4(3,2218,418);
  `device_slave_connections_TB_CONFIG_4(3,2219,419);
  `device_slave_connections_TB_CONFIG_4(3,2220,420);
  `device_slave_connections_TB_CONFIG_4(3,2221,421);
  `device_slave_connections_TB_CONFIG_4(3,2222,422);
  `device_slave_connections_TB_CONFIG_4(3,2223,423);
  `device_slave_connections_TB_CONFIG_4(3,2224,424);
  `device_slave_connections_TB_CONFIG_4(3,2225,425);
  `device_slave_connections_TB_CONFIG_4(3,2226,426);
  `device_slave_connections_TB_CONFIG_4(3,2227,427);
  `device_slave_connections_TB_CONFIG_4(3,2228,428);
  `device_slave_connections_TB_CONFIG_4(3,2229,429);
  `device_slave_connections_TB_CONFIG_4(3,2230,430);
  `device_slave_connections_TB_CONFIG_4(3,2231,431);
  `device_slave_connections_TB_CONFIG_4(3,2232,432);
  `device_slave_connections_TB_CONFIG_4(3,2233,433);
  `device_slave_connections_TB_CONFIG_4(3,2234,434);
  `device_slave_connections_TB_CONFIG_4(3,2235,435);
  `device_slave_connections_TB_CONFIG_4(3,2236,436);
  `device_slave_connections_TB_CONFIG_4(3,2237,437);
  `device_slave_connections_TB_CONFIG_4(3,2238,438);
  `device_slave_connections_TB_CONFIG_4(3,2239,439);
  `device_slave_connections_TB_CONFIG_4(3,2240,440);
  `device_slave_connections_TB_CONFIG_4(3,2241,441);
  `device_slave_connections_TB_CONFIG_4(3,2242,442);
  `device_slave_connections_TB_CONFIG_4(3,2243,443);
  `device_slave_connections_TB_CONFIG_4(3,2244,444);
  `device_slave_connections_TB_CONFIG_4(3,2245,445);
  `device_slave_connections_TB_CONFIG_4(3,2246,446);
  `device_slave_connections_TB_CONFIG_4(3,2247,447);
  `device_slave_connections_TB_CONFIG_4(3,2248,448);
  `device_slave_connections_TB_CONFIG_4(3,2249,449);
	*/
	
  `elsif TB_CONFIG_2
  `device_slave_connections_N(16,0);
  `device_slave_connections_N(17,1);
  `device_slave_connections_N(18,2);
  `device_slave_connections_N(19,3);
  `device_slave_connections_N(20,4);
  `device_slave_connections_N(21,5);
  `device_slave_connections_N(22,6);
  `device_slave_connections_N(23,7);

	`elsif TB_CONFIG_3
  `device_slave_connections_N(16,0);
  `device_slave_connections_N(17,1);
  `device_slave_connections_N(18,2);
  `device_slave_connections_N(19,3);
  `device_slave_connections_N(20,4);
  `device_slave_connections_N(21,5);
  `device_slave_connections_N(22,6);
  `device_slave_connections_N(23,7);
  `device_slave_connections_N(24,8);
  `device_slave_connections_N(25,9);
  `device_slave_connections_N(26,10);
  `device_slave_connections_N(27,11);
  `device_slave_connections_N(28,12);
  `device_slave_connections_N(29,13);
  `device_slave_connections_N(30,14);
  `device_slave_connections_N(31,15);
	`endif

  //=======================
  // Mux --> Host 
  //=======================
  force axis_if_H.slave_if[0].tvalid        =   `TOP.mx2ho_tx_port.tvalid;      
  force axis_if_H.slave_if[0].tlast         =   `TOP.mx2ho_tx_port.tlast;              
  force axis_if_H.slave_if[0].tuser         =   `TOP.mx2ho_tx_port.tuser_vendor;                
  force axis_if_H.slave_if[0].tdata         =   `TOP.mx2ho_tx_port.tdata;                
  force axis_if_H.slave_if[0].tkeep         =   `TOP.mx2ho_tx_port.tkeep; 
  force axis_if_H.slave_if[0].tready        =   `TOP.mx2ho_tx_port.tready;
  
  //===============================================================================
  //Added just to remove the assertion error : Offending '(!$isunknown(tvalid/tready))'
  //===============================================================================
       force top_tb.mx2fn_rx_remap[0].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[2].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[3].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[4].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[5].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[6].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[7].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[8].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[9].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[10].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[11].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[12].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[13].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[14].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[15].tready = 1'b1;
      `ifdef TB_CONFIG_4
       force top_tb.mx2fn_rx_remap[16].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[17].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[18].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[19].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[20].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[21].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[22].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[23].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[24].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[25].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[26].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[27].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[28].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[29].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[30].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[31].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[32].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[33].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[34].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[35].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[36].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[37].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[38].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[39].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[40].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[41].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[42].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[43].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[44].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[45].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[46].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[47].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[48].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[49].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[50].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[51].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[52].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[53].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[54].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[55].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[56].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[57].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[58].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[59].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[60].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[61].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[62].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[63].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[64].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[65].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[66].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[67].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[68].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[69].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[70].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[71].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[72].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[73].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[74].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[75].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[76].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[77].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[78].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[79].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[80].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[81].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[82].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[83].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[84].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[85].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[86].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[87].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[88].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[89].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[90].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[91].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[92].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[93].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[94].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[95].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[96].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[97].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[98].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[99].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[100].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[101].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[102].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[103].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[104].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[105].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[106].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[107].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[108].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[109].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[110].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[111].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[112].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[113].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[114].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[115].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[116].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[117].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[118].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[119].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[120].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[121].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[122].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[123].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[124].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[125].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[126].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[127].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[128].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[129].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[130].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[131].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[132].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[133].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[134].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[135].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[136].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[137].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[138].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[139].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[140].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[141].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[142].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[143].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[144].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[145].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[146].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[147].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[148].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[149].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[150].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[151].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[152].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[153].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[154].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[155].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[156].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[157].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[158].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[159].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[160].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[161].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[162].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[163].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[164].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[165].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[166].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[167].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[168].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[169].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[170].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[171].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[172].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[173].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[174].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[175].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[176].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[177].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[178].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[179].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[180].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[181].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[182].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[183].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[184].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[185].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[186].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[187].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[188].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[189].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[190].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[191].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[192].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[193].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[194].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[195].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[196].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[197].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[198].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[199].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[200].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[201].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[202].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[203].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[204].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[205].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[206].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[207].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[208].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[209].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[210].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[211].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[212].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[213].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[214].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[215].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[216].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[217].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[218].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[219].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[220].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[221].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[222].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[223].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[224].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[225].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[226].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[227].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[228].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[229].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[230].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[231].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[232].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[233].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[234].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[235].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[236].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[237].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[238].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[239].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[240].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[241].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[242].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[243].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[244].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[245].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[246].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[247].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[248].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[249].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[250].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[251].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[252].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[253].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[254].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[255].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[256].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[257].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[258].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[259].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[260].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[261].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[262].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[263].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[264].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[265].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[266].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[267].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[268].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[269].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[270].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[271].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[272].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[273].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[274].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[275].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[276].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[277].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[278].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[279].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[280].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[281].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[282].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[283].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[284].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[285].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[286].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[287].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[288].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[289].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[290].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[291].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[292].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[293].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[294].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[295].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[296].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[297].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[298].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[299].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[300].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[301].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[302].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[303].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[304].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[305].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[306].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[307].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[308].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[309].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[310].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[311].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[312].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[313].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[314].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[315].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[316].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[317].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[318].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[319].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[320].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[321].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[322].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[323].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[324].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[325].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[326].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[327].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[328].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[329].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[330].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[331].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[332].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[333].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[334].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[335].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[336].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[337].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[338].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[339].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[340].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[341].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[342].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[343].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[344].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[345].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[346].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[347].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[348].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[349].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[350].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[351].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[352].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[353].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[354].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[355].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[356].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[357].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[358].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[359].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[360].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[361].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[362].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[363].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[364].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[365].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[366].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[367].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[368].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[369].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[370].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[371].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[372].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[373].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[374].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[375].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[376].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[377].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[378].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[379].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[380].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[381].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[382].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[383].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[384].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[385].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[386].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[387].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[388].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[389].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[390].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[391].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[392].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[393].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[394].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[395].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[396].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[397].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[398].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[399].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[400].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[401].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[402].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[403].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[404].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[405].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[406].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[407].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[408].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[409].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[410].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[411].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[412].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[413].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[414].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[415].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[416].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[417].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[418].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[419].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[420].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[421].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[422].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[423].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[424].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[425].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[426].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[427].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[428].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[429].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[430].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[431].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[432].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[433].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[434].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[435].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[436].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[437].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[438].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[439].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[440].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[441].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[442].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[443].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[444].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[445].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[446].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[447].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[448].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[449].tready = 1'b1;
			 force top_tb.mx2fn_rx_remap[450].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[451].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[452].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[453].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[454].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[455].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[456].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[457].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[458].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[459].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[460].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[461].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[462].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[463].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[464].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[465].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[466].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[467].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[468].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[469].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[470].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[471].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[472].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[473].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[474].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[475].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[476].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[477].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[478].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[479].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[480].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[481].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[482].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[483].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[484].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[485].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[486].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[487].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[488].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[489].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[490].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[491].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[492].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[493].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[494].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[495].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[496].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[497].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[498].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[499].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[500].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[501].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[502].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[503].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[504].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[505].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[506].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[507].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[508].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[509].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[510].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[511].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[512].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[513].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[514].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[515].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[516].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[517].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[518].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[519].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[520].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[521].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[522].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[523].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[524].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[525].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[526].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[527].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[528].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[529].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[530].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[531].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[532].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[533].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[534].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[535].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[536].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[537].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[538].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[539].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[540].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[541].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[542].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[543].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[544].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[545].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[546].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[547].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[548].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[549].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[550].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[551].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[552].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[553].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[554].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[555].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[556].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[557].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[558].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[559].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[560].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[561].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[562].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[563].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[564].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[565].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[566].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[567].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[568].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[569].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[570].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[571].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[572].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[573].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[574].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[575].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[576].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[577].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[578].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[579].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[580].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[581].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[582].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[583].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[584].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[585].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[586].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[587].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[588].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[589].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[590].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[591].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[592].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[593].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[594].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[595].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[596].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[597].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[598].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[599].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[600].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[601].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[602].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[603].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[604].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[605].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[606].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[607].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[608].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[609].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[610].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[611].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[612].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[613].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[614].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[615].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[616].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[617].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[618].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[619].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[620].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[621].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[622].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[623].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[624].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[625].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[626].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[627].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[628].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[629].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[630].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[631].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[632].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[633].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[634].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[635].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[636].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[637].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[638].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[639].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[640].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[641].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[642].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[643].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[644].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[645].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[646].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[647].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[648].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[649].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[650].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[651].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[652].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[653].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[654].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[655].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[656].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[657].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[658].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[659].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[660].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[661].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[662].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[663].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[664].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[665].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[666].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[667].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[668].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[669].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[670].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[671].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[672].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[673].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[674].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[675].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[676].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[677].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[678].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[679].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[680].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[681].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[682].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[683].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[684].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[685].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[686].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[687].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[688].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[689].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[690].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[691].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[692].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[693].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[694].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[695].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[696].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[697].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[698].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[699].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[700].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[701].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[702].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[703].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[704].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[705].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[706].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[707].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[708].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[709].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[710].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[711].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[712].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[713].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[714].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[715].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[716].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[717].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[718].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[719].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[720].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[721].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[722].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[723].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[724].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[725].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[726].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[727].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[728].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[729].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[730].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[731].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[732].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[733].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[734].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[735].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[736].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[737].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[738].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[739].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[740].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[741].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[742].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[743].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[744].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[745].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[746].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[747].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[748].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[749].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[750].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[751].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[752].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[753].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[754].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[755].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[756].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[757].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[758].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[759].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[760].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[761].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[762].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[763].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[764].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[765].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[766].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[767].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[768].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[769].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[770].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[771].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[772].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[773].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[774].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[775].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[776].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[777].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[778].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[779].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[780].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[781].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[782].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[783].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[784].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[785].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[786].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[787].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[788].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[789].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[790].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[791].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[792].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[793].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[794].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[795].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[796].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[797].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[798].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[799].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[800].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[801].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[802].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[803].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[804].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[805].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[806].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[807].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[808].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[809].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[810].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[811].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[812].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[813].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[814].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[815].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[816].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[817].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[818].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[819].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[820].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[821].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[822].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[823].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[824].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[825].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[826].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[827].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[828].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[829].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[830].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[831].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[832].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[833].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[834].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[835].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[836].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[837].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[838].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[839].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[840].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[841].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[842].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[843].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[844].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[845].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[846].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[847].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[848].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[849].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[850].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[851].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[852].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[853].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[854].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[855].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[856].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[857].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[858].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[859].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[860].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[861].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[862].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[863].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[864].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[865].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[866].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[867].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[868].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[869].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[870].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[871].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[872].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[873].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[874].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[875].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[876].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[877].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[878].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[879].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[880].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[881].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[882].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[883].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[884].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[885].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[886].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[887].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[888].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[889].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[890].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[891].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[892].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[893].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[894].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[895].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[896].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[897].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[898].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[899].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[900].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[901].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[902].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[903].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[904].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[905].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[906].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[907].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[908].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[909].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[910].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[911].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[912].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[913].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[914].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[915].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[916].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[917].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[918].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[919].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[920].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[921].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[922].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[923].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[924].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[925].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[926].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[927].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[928].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[929].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[930].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[931].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[932].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[933].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[934].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[935].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[936].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[937].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[938].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[939].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[940].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[941].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[942].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[943].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[944].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[945].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[946].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[947].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[948].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[949].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[950].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[951].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[952].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[953].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[954].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[955].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[956].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[957].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[958].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[959].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[960].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[961].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[962].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[963].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[964].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[965].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[966].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[967].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[968].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[969].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[970].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[971].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[972].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[973].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[974].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[975].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[976].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[977].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[978].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[979].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[980].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[981].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[982].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[983].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[984].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[985].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[986].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[987].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[988].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[989].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[990].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[991].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[992].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[993].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[994].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[995].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[996].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[997].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[998].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[999].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1000].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1001].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1002].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1003].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1004].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1005].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1006].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1007].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1008].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1009].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1010].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1011].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1012].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1013].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1014].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1015].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1016].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1017].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1018].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1019].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1020].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1021].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1022].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1023].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1024].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1025].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1026].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1027].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1028].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1029].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1030].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1031].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1032].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1033].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1034].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1035].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1036].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1037].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1038].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1039].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1040].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1041].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1042].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1043].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1044].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1045].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1046].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1047].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1048].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1049].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1050].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1051].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1052].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1053].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1054].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1055].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1056].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1057].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1058].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1059].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1060].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1061].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1062].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1063].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1064].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1065].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1066].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1067].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1068].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1069].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1070].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1071].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1072].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1073].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1074].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1075].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1076].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1077].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1078].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1079].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1080].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1081].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1082].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1083].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1084].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1085].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1086].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1087].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1088].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1089].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1090].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1091].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1092].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1093].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1094].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1095].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1096].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1097].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1098].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1099].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1100].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1101].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1102].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1103].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1104].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1105].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1106].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1107].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1108].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1109].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1110].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1111].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1112].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1113].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1114].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1115].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1116].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1117].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1118].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1119].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1120].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1121].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1122].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1123].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1124].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1125].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1126].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1127].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1128].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1129].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1130].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1131].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1132].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1133].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1134].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1135].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1136].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1137].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1138].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1139].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1140].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1141].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1142].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1143].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1144].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1145].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1146].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1147].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1148].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1149].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1150].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1151].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1152].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1153].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1154].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1155].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1156].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1157].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1158].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1159].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1160].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1161].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1162].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1163].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1164].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1165].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1166].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1167].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1168].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1169].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1170].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1171].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1172].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1173].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1174].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1175].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1176].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1177].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1178].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1179].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1180].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1181].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1182].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1183].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1184].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1185].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1186].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1187].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1188].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1189].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1190].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1191].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1192].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1193].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1194].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1195].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1196].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1197].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1198].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1199].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1200].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1201].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1202].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1203].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1204].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1205].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1206].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1207].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1208].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1209].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1210].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1211].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1212].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1213].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1214].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1215].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1216].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1217].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1218].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1219].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1220].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1221].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1222].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1223].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1224].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1225].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1226].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1227].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1228].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1229].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1230].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1231].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1232].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1233].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1234].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1235].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1236].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1237].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1238].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1239].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1240].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1241].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1242].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1243].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1244].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1245].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1246].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1247].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1248].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1249].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1250].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1251].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1252].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1253].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1254].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1255].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1256].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1257].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1258].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1259].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1260].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1261].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1262].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1263].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1264].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1265].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1266].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1267].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1268].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1269].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1270].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1271].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1272].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1273].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1274].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1275].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1276].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1277].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1278].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1279].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1280].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1281].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1282].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1283].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1284].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1285].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1286].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1287].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1288].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1289].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1290].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1291].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1292].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1293].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1294].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1295].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1296].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1297].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1298].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1299].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1300].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1301].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1302].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1303].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1304].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1305].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1306].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1307].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1308].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1309].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1310].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1311].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1312].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1313].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1314].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1315].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1316].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1317].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1318].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1319].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1320].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1321].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1322].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1323].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1324].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1325].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1326].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1327].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1328].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1329].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1330].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1331].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1332].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1333].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1334].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1335].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1336].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1337].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1338].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1339].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1340].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1341].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1342].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1343].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1344].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1345].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1346].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1347].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1348].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1349].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1350].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1351].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1352].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1353].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1354].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1355].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1356].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1357].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1358].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1359].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1360].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1361].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1362].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1363].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1364].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1365].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1366].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1367].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1368].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1369].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1370].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1371].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1372].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1373].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1374].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1375].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1376].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1377].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1378].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1379].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1380].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1381].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1382].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1383].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1384].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1385].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1386].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1387].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1388].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1389].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1390].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1391].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1392].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1393].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1394].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1395].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1396].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1397].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1398].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1399].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1400].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1401].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1402].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1403].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1404].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1405].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1406].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1407].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1408].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1409].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1410].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1411].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1412].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1413].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1414].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1415].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1416].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1417].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1418].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1419].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1420].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1421].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1422].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1423].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1424].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1425].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1426].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1427].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1428].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1429].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1430].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1431].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1432].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1433].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1434].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1435].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1436].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1437].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1438].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1439].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1440].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1441].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1442].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1443].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1444].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1445].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1446].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1447].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1448].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1449].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1450].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1451].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1452].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1453].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1454].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1455].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1456].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1457].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1458].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1459].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1460].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1461].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1462].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1463].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1464].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1465].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1466].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1467].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1468].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1469].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1470].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1471].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1472].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1473].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1474].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1475].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1476].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1477].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1478].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1479].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1480].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1481].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1482].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1483].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1484].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1485].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1486].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1487].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1488].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1489].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1490].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1491].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1492].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1493].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1494].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1495].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1496].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1497].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1498].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1499].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1500].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1501].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1502].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1503].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1504].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1505].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1506].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1507].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1508].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1509].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1510].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1511].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1512].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1513].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1514].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1515].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1516].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1517].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1518].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1519].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1520].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1521].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1522].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1523].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1524].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1525].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1526].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1527].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1528].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1529].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1530].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1531].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1532].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1533].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1534].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1535].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1536].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1537].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1538].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1539].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1540].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1541].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1542].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1543].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1544].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1545].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1546].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1547].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1548].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1549].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1550].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1551].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1552].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1553].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1554].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1555].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1556].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1557].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1558].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1559].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1560].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1561].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1562].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1563].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1564].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1565].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1566].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1567].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1568].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1569].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1570].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1571].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1572].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1573].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1574].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1575].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1576].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1577].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1578].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1579].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1580].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1581].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1582].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1583].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1584].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1585].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1586].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1587].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1588].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1589].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1590].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1591].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1592].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1593].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1594].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1595].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1596].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1597].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1598].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1599].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1600].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1601].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1602].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1603].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1604].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1605].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1606].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1607].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1608].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1609].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1610].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1611].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1612].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1613].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1614].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1615].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1616].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1617].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1618].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1619].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1620].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1621].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1622].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1623].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1624].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1625].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1626].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1627].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1628].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1629].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1630].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1631].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1632].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1633].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1634].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1635].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1636].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1637].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1638].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1639].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1640].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1641].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1642].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1643].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1644].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1645].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1646].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1647].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1648].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1649].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1650].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1651].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1652].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1653].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1654].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1655].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1656].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1657].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1658].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1659].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1660].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1661].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1662].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1663].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1664].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1665].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1666].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1667].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1668].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1669].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1670].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1671].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1672].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1673].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1674].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1675].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1676].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1677].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1678].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1679].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1680].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1681].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1682].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1683].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1684].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1685].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1686].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1687].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1688].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1689].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1690].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1691].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1692].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1693].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1694].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1695].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1696].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1697].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1698].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1699].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1700].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1701].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1702].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1703].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1704].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1705].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1706].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1707].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1708].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1709].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1710].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1711].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1712].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1713].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1714].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1715].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1716].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1717].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1718].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1719].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1720].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1721].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1722].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1723].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1724].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1725].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1726].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1727].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1728].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1729].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1730].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1731].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1732].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1733].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1734].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1735].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1736].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1737].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1738].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1739].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1740].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1741].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1742].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1743].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1744].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1745].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1746].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1747].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1748].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1749].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1750].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1751].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1752].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1753].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1754].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1755].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1756].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1757].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1758].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1759].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1760].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1761].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1762].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1763].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1764].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1765].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1766].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1767].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1768].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1769].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1770].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1771].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1772].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1773].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1774].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1775].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1776].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1777].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1778].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1779].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1780].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1781].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1782].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1783].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1784].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1785].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1786].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1787].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1788].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1789].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1790].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1791].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1792].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1793].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1794].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1795].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1796].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1797].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1798].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1799].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1800].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1801].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1802].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1803].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1804].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1805].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1806].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1807].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1808].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1809].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1810].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1811].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1812].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1813].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1814].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1815].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1816].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1817].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1818].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1819].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1820].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1821].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1822].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1823].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1824].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1825].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1826].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1827].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1828].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1829].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1830].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1831].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1832].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1833].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1834].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1835].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1836].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1837].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1838].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1839].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1840].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1841].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1842].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1843].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1844].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1845].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1846].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1847].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1848].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1849].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1850].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1851].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1852].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1853].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1854].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1855].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1856].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1857].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1858].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1859].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1860].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1861].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1862].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1863].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1864].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1865].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1866].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1867].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1868].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1869].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1870].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1871].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1872].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1873].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1874].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1875].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1876].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1877].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1878].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1879].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1880].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1881].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1882].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1883].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1884].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1885].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1886].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1887].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1888].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1889].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1890].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1891].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1892].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1893].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1894].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1895].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1896].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1897].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1898].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1899].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1900].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1901].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1902].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1903].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1904].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1905].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1906].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1907].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1908].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1909].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1910].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1911].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1912].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1913].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1914].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1915].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1916].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1917].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1918].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1919].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1920].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1921].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1922].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1923].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1924].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1925].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1926].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1927].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1928].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1929].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1930].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1931].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1932].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1933].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1934].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1935].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1936].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1937].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1938].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1939].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1940].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1941].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1942].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1943].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1944].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1945].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1946].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1947].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1948].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1949].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1950].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1951].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1952].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1953].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1954].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1955].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1956].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1957].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1958].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1959].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1960].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1961].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1962].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1963].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1964].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1965].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1966].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1967].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1968].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1969].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1970].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1971].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1972].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1973].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1974].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1975].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1976].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1977].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1978].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1979].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1980].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1981].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1982].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1983].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1984].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1985].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1986].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1987].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1988].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1989].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1990].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1991].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1992].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1993].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1994].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1995].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1996].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1997].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1998].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[1999].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[2000].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[2001].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[2002].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[2003].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[2004].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[2005].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[2006].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[2007].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[2008].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[2009].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[2010].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[2011].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[2012].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[2013].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[2014].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[2015].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[2016].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[2017].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[2018].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[2019].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[2020].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[2021].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[2022].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[2023].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[2024].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[2025].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[2026].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[2027].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[2028].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[2029].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[2030].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[2031].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[2032].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[2033].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[2034].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[2035].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[2036].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[2037].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[2038].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[2039].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[2040].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[2041].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[2042].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[2043].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[2044].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[2045].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[2046].tready = 1'b1;
       force top_tb.mx2fn_rx_remap[2047].tready = 1'b1;

		`elsif TB_CONFIG_2
    force top_tb.mx2fn_rx_remap[16].tready = 1'b1;
    force top_tb.mx2fn_rx_remap[17].tready = 1'b1;
    force top_tb.mx2fn_rx_remap[18].tready = 1'b1;
    force top_tb.mx2fn_rx_remap[19].tready = 1'b1;
    force top_tb.mx2fn_rx_remap[20].tready = 1'b1;
    force top_tb.mx2fn_rx_remap[21].tready = 1'b1;
    force top_tb.mx2fn_rx_remap[22].tready = 1'b1;
    force top_tb.mx2fn_rx_remap[23].tready = 1'b1;
    
		`elsif TB_CONFIG_3
    force top_tb.mx2fn_rx_remap[16].tready = 1'b1;
    force top_tb.mx2fn_rx_remap[17].tready = 1'b1;
    force top_tb.mx2fn_rx_remap[18].tready = 1'b1;
    force top_tb.mx2fn_rx_remap[19].tready = 1'b1;
    force top_tb.mx2fn_rx_remap[20].tready = 1'b1;
    force top_tb.mx2fn_rx_remap[21].tready = 1'b1;
    force top_tb.mx2fn_rx_remap[22].tready = 1'b1;
    force top_tb.mx2fn_rx_remap[23].tready = 1'b1;
    force top_tb.mx2fn_rx_remap[24].tready = 1'b1;
    force top_tb.mx2fn_rx_remap[25].tready = 1'b1;
    force top_tb.mx2fn_rx_remap[26].tready = 1'b1;
    force top_tb.mx2fn_rx_remap[27].tready = 1'b1;
    force top_tb.mx2fn_rx_remap[28].tready = 1'b1;
    force top_tb.mx2fn_rx_remap[29].tready = 1'b1;
    force top_tb.mx2fn_rx_remap[30].tready = 1'b1;
    force top_tb.mx2fn_rx_remap[31].tready = 1'b1;
		`endif

    `ifdef TB_CONFIG_4   //We are not using below mentioned ports from 248 to 449 for last VIP
      force TB4_axis_if_D3.slave_if[248].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[249].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[250].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[251].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[252].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[253].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[254].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[255].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[256].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[257].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[258].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[259].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[260].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[261].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[262].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[263].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[264].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[265].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[266].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[267].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[268].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[269].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[270].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[271].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[272].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[273].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[274].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[275].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[276].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[277].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[278].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[279].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[280].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[281].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[282].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[283].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[284].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[285].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[286].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[287].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[288].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[289].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[290].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[291].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[292].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[293].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[294].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[295].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[296].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[297].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[298].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[299].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[300].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[301].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[302].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[303].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[304].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[305].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[306].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[307].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[308].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[309].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[310].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[311].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[312].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[313].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[314].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[315].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[316].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[317].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[318].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[319].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[320].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[321].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[322].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[323].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[324].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[325].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[326].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[327].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[328].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[329].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[330].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[331].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[332].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[333].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[334].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[335].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[336].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[337].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[338].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[339].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[340].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[341].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[342].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[343].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[344].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[345].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[346].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[347].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[348].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[349].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[350].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[351].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[352].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[353].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[354].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[355].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[356].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[357].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[358].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[359].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[360].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[361].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[362].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[363].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[364].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[365].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[366].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[367].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[368].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[369].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[370].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[371].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[372].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[373].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[374].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[375].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[376].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[377].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[378].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[379].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[380].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[381].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[382].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[383].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[384].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[385].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[386].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[387].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[388].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[389].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[390].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[391].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[392].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[393].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[394].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[395].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[396].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[397].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[398].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[399].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[400].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[401].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[402].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[403].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[404].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[405].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[406].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[407].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[408].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[409].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[410].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[411].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[412].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[413].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[414].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[415].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[416].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[417].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[418].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[419].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[420].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[421].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[422].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[423].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[424].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[425].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[426].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[427].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[428].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[429].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[430].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[431].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[432].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[433].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[434].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[435].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[436].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[437].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[438].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[439].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[440].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[441].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[442].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[443].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[444].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[445].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[446].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[447].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[448].tvalid = 1'b0 ;
      force TB4_axis_if_D3.slave_if[449].tvalid = 1'b0 ;
     `endif
end

always @(posedge top_tb.clk)
  if(top_tb.rst_n)
    begin
      top_tb.mx2ho_tx_remap.tready <= 1'b1;
    end

endmodule
