// Copyright (C) 2023 Intel Corporation
// SPDX-License-Identifier: MIT

`define toggle_tready(PORT) \
 begin\
  if(i<=(no_of_transactions/3))\    
    force top_tb.pf_vf_mux_a.mx2fn_rx_port[``PORT``].tready         =  1;\
  else if ((i>=(no_of_transactions/3)) && (i<=(2*no_of_transactions/3)))\
    force top_tb.pf_vf_mux_a.mx2fn_rx_port[``PORT``].tready         =  0;\ 
  else\ 
    force top_tb.pf_vf_mux_a.mx2fn_rx_port[``PORT``].tready         =  1;\ 
 end\

`define fifo_error_check(PORT)\
begin\
 if(top_tb.pf_vf_mux_a.switch.N_mux[``PORT``].out_q.fifo_cntr == 2)\ 
   begin\
    `uvm_info("body", "OVERFLOW_FIFO_ERR_``PORT``", UVM_LOW)\
     force top_tb.pf_vf_mux_a.switch.N_mux[``PORT``].out_q.fifo_wen = 1;\
     @(posedge top_tb.pf_vf_mux_a.switch.N_mux[``PORT``].out_q.clk);\
     release top_tb.pf_vf_mux_a.switch.N_mux[``PORT``].out_q.fifo_wen;\
   end\ 
 if(i == 0)\
   begin\
    `uvm_info("body", "UNDERFLOW_FIFO_ERR_``PORT``", UVM_LOW)\
     force top_tb.pf_vf_mux_a.switch.N_mux[``PORT``].out_q.fifo_ren = 1;\
     @(posedge top_tb.pf_vf_mux_a.switch.N_mux[``PORT``].out_q.clk);\
     release top_tb.pf_vf_mux_a.switch.N_mux[``PORT``].out_q.fifo_ren;\
     @(posedge top_tb.pf_vf_mux_a.switch.N_mux[``PORT``].out_q.clk);\
     force top_tb.pf_vf_mux_a.switch.N_mux[``PORT``].out_q.fifo_ren = 1;\
     @(posedge top_tb.pf_vf_mux_a.switch.N_mux[``PORT``].out_q.clk);\
     release top_tb.pf_vf_mux_a.switch.N_mux[``PORT``].out_q.fifo_ren;\
     @(posedge top_tb.pf_vf_mux_a.switch.N_mux[``PORT``].out_q.clk);\
     force top_tb.pf_vf_mux_a.switch.N_mux[``PORT``].out_q.fifo_ren = 1;\
     @(posedge top_tb.pf_vf_mux_a.switch.N_mux[``PORT``].out_q.clk);\
     release top_tb.pf_vf_mux_a.switch.N_mux[``PORT``].out_q.fifo_ren;\
   end\
end\  

class pf_vf_mux_master_fifo_error_seq extends uvm_sequence;
    
     rand bit local_vf_active       ;
     rand bit [2:0] local_pf_num    ;
     rand bit [10:0] local_vf_num   ;
     bit [9:0] local_tlp_length;
     bit [255:0] local_payload , random_value, local_my_payload;
     rand int no_of_transactions ;
     
    `ifdef TB_CONFIG_4
     bit vf_active_array[1] ;
     bit[10:0] vf_num_array[1];
     `elsif TB_CONFIG_3
     bit vf_active_array[4] ;
     bit[10:0] vf_num_array[4];
     `elsif TB_CONFIG_2
     bit vf_active_array[3] ;
     bit[10:0] vf_num_array[3];
     `else 
     bit vf_active_array[2] ;
     bit[10:0] vf_num_array[2];
     `endif

     int vf_va = 0;
     int count;

    `uvm_object_utils(pf_vf_mux_master_fifo_error_seq);

  /** Declare a typed sequencer object that the sequence can access */
  `uvm_declare_p_sequencer(pf_vf_mux_virtual_sequencer)


    function new (string name = "pf_vf_mux_master_fifo_error_seq");
        super.new(name);
    endfunction : new

     virtual function void build_phase(uvm_phase phase);
        `uvm_info ("build_phase", "Entered PF0 Traffic Sequence Build Phase...",UVM_LOW);
      endfunction: build_phase


    task body();
        pf_vf_mux_request_sequence master_seq;

        super.body(); 
      	`uvm_info(get_name(), "Entering PF0 Traffic sequence...", UVM_LOW)
        `uvm_info(get_name(), "Starting master sequence on Host master sequencer", UVM_LOW)

        `ifdef TB_CONFIG_4 
        vf_active_array = '{'h1};
        vf_num_array    = '{'h0};
        vf_va = 1;
        `elsif TB_CONFIG_3 
        vf_active_array = '{'h0,'h1,'h1,'h1};
        vf_num_array    = '{'h0,'h0,'h7ff,`RANDOM_VF};
        vf_va = 4;
        `elsif TB_CONFIG_2 
        vf_active_array = '{'h0,'h1,'h1};
        vf_num_array    = '{'h0,'h0,'h7ff};
        vf_va = 3;
        `else 
        vf_active_array = '{'h0,'h1};
        vf_num_array    = '{'h0,'h0};
        vf_va = 2;
        `endif

          for(int k = 0; k < vf_va; k++) begin //{
         `ifdef TB_CONFIG_4
          for(int t = 0; t < 2048; t++) begin //{
         `else
          for(int j = 0; j < 8; j++) begin //{
         `endif
          for(int i = 0; i < no_of_transactions; i++) begin
            //===============================================
            // Generating the payload w.r.t TLP length field
            //===============================================
            local_vf_active = vf_active_array[k];
           `ifdef TB_CONFIG_4
            local_pf_num = 0;
            local_vf_num = t;
           `else
            local_pf_num = j;
            local_vf_num = vf_num_array[k];
           `endif
            local_tlp_length = $urandom_range(1,64) ;
            local_payload = 'h0;
            local_my_payload = 'h0;
            assert(std::randomize(random_value));      
            `uvm_info("body", $sformatf("LOCAL_PF_NUM = %d and LOCAL_VF_NUM = %d and LOCAL_VF_ACTIVE = %d",local_pf_num,local_vf_num,local_vf_active), UVM_LOW)
            for(int l=0; l < (local_tlp_length*32); l++) local_my_payload[l] = 1'b1;
            local_payload = (random_value) & local_my_payload;
            `uvm_info("body", $sformatf("TLP Length = %h and Payload = %h and Random Value generated = %h",local_tlp_length,local_payload,random_value), UVM_LOW)

              `ifdef TB_CONFIG_1
              if (local_pf_num==0 && local_vf_num==0 && local_vf_active==0)
               `fifo_error_check(0)              
              else if (local_pf_num==1 && local_vf_num==0 && local_vf_active==0) 
                `fifo_error_check(1)                   
              else if (local_pf_num==2 && local_vf_num==0 && local_vf_active==0) 
                 `fifo_error_check(2)                  
              else if (local_pf_num==3 && local_vf_num==0 && local_vf_active==0) 
                  `fifo_error_check(3)                 
              else if (local_pf_num==4 && local_vf_num==0 && local_vf_active==0) 
                  `fifo_error_check(4)                                         
              else if (local_pf_num==5 && local_vf_num==0 && local_vf_active==0) 
                   `fifo_error_check(5)                                        
              else if (local_pf_num==6 && local_vf_num==0 && local_vf_active==0) 
                   `fifo_error_check(6)                         
              else if (local_pf_num==7 && local_vf_num==0 && local_vf_active==0) 
                    `fifo_error_check(7)                                       
              else if (local_pf_num==0 && local_vf_num==0 && local_vf_active==1) 
                    `fifo_error_check(8)                                       
              else if (local_pf_num==1 && local_vf_num==0 && local_vf_active==1) 
                    `fifo_error_check(9)     
              else if (local_pf_num==2 && local_vf_num==0 && local_vf_active==1) 
                   `fifo_error_check(10)                    
              else if (local_pf_num==3 && local_vf_num==0 && local_vf_active==1) 
                   `fifo_error_check(11)                    
              else if (local_pf_num==4 && local_vf_num==0 && local_vf_active==1) 
                   `fifo_error_check(12)     
              else if (local_pf_num==5 && local_vf_num==0 && local_vf_active==1) 
                   `fifo_error_check(13)                    
              else if (local_pf_num==6 && local_vf_num==0 && local_vf_active==1) 
                   `fifo_error_check(14)                    
              else if (local_pf_num==7 && local_vf_num==0 && local_vf_active==1) 
                   `fifo_error_check(15)

              `elsif TB_CONFIG_2
              if (local_pf_num==0 && local_vf_num==0 && local_vf_active==0)
               `fifo_error_check(0)              
              else if (local_pf_num==1 && local_vf_num==0 && local_vf_active==0) 
                `fifo_error_check(1)                   
              else if (local_pf_num==2 && local_vf_num==0 && local_vf_active==0) 
                 `fifo_error_check(2)                  
              else if (local_pf_num==3 && local_vf_num==0 && local_vf_active==0) 
                  `fifo_error_check(3)                 
              else if (local_pf_num==4 && local_vf_num==0 && local_vf_active==0) 
                  `fifo_error_check(4)                                         
              else if (local_pf_num==5 && local_vf_num==0 && local_vf_active==0) 
                   `fifo_error_check(5)                                        
              else if (local_pf_num==6 && local_vf_num==0 && local_vf_active==0) 
                   `fifo_error_check(6)                         
              else if (local_pf_num==7 && local_vf_num==0 && local_vf_active==0) 
                    `fifo_error_check(7)                                       
              else if (local_pf_num==0 && local_vf_num==0 && local_vf_active==1) 
                    `fifo_error_check(8)                                       
              else if (local_pf_num==1 && local_vf_num==0 && local_vf_active==1) 
                    `fifo_error_check(9)     
              else if (local_pf_num==2 && local_vf_num==0 && local_vf_active==1) 
                   `fifo_error_check(10)                    
              else if (local_pf_num==3 && local_vf_num==0 && local_vf_active==1) 
                   `fifo_error_check(11)                    
              else if (local_pf_num==4 && local_vf_num==0 && local_vf_active==1) 
                   `fifo_error_check(12)     
              else if (local_pf_num==5 && local_vf_num==0 && local_vf_active==1) 
                   `fifo_error_check(13)                    
              else if (local_pf_num==6 && local_vf_num==0 && local_vf_active==1) 
                   `fifo_error_check(14)                    
              else if (local_pf_num==7 && local_vf_num==0 && local_vf_active==1) 
                    `fifo_error_check(15)
              else if (local_pf_num==0 && local_vf_num=='h7ff && local_vf_active==1) 
                    `fifo_error_check(16)                                           
              else if (local_pf_num==1 && local_vf_num=='h7ff && local_vf_active==1) 
                    `fifo_error_check(17)                                           
              else if (local_pf_num==2 && local_vf_num=='h7ff && local_vf_active==1) 
                   `fifo_error_check(18)                                            
              else if (local_pf_num==3 && local_vf_num=='h7ff && local_vf_active==1) 
                   `fifo_error_check(19)                                            
              else if (local_pf_num==4 && local_vf_num=='h7ff && local_vf_active==1) 
                   `fifo_error_check(20)                                           
              else if (local_pf_num==5 && local_vf_num=='h7ff && local_vf_active==1) 
                   `fifo_error_check(21)                                        
              else if (local_pf_num==6 && local_vf_num=='h7ff && local_vf_active==1) 
                   `fifo_error_check(22)                                            
              else if (local_pf_num==7 && local_vf_num=='h7ff && local_vf_active==1) 
                    `fifo_error_check(23)

              `elsif TB_CONFIG_3
              if (local_pf_num==0 && local_vf_num==0 && local_vf_active==0)
               `fifo_error_check(0)              
              else if (local_pf_num==1 && local_vf_num==0 && local_vf_active==0) 
                `fifo_error_check(1)                   
              else if (local_pf_num==2 && local_vf_num==0 && local_vf_active==0) 
                 `fifo_error_check(2)                  
              else if (local_pf_num==3 && local_vf_num==0 && local_vf_active==0) 
                  `fifo_error_check(3)                 
              else if (local_pf_num==4 && local_vf_num==0 && local_vf_active==0) 
                  `fifo_error_check(4)                                         
              else if (local_pf_num==5 && local_vf_num==0 && local_vf_active==0) 
                   `fifo_error_check(5)                                        
              else if (local_pf_num==6 && local_vf_num==0 && local_vf_active==0) 
                   `fifo_error_check(6)                         
              else if (local_pf_num==7 && local_vf_num==0 && local_vf_active==0) 
                    `fifo_error_check(7)                                       
              else if (local_pf_num==0 && local_vf_num==0 && local_vf_active==1) 
                    `fifo_error_check(8)                                       
              else if (local_pf_num==1 && local_vf_num==0 && local_vf_active==1) 
                    `fifo_error_check(9)     
              else if (local_pf_num==2 && local_vf_num==0 && local_vf_active==1) 
                   `fifo_error_check(10)                    
              else if (local_pf_num==3 && local_vf_num==0 && local_vf_active==1) 
                   `fifo_error_check(11)                    
              else if (local_pf_num==4 && local_vf_num==0 && local_vf_active==1) 
                   `fifo_error_check(12)     
              else if (local_pf_num==5 && local_vf_num==0 && local_vf_active==1) 
                   `fifo_error_check(13)                    
              else if (local_pf_num==6 && local_vf_num==0 && local_vf_active==1) 
                   `fifo_error_check(14)                    
              else if (local_pf_num==7 && local_vf_num==0 && local_vf_active==1) 
                    `fifo_error_check(15)
              else if (local_pf_num==0 && local_vf_num=='h7ff && local_vf_active==1) 
                    `fifo_error_check(16)                                           
              else if (local_pf_num==1 && local_vf_num=='h7ff && local_vf_active==1) 
                    `fifo_error_check(17)                                           
              else if (local_pf_num==2 && local_vf_num=='h7ff && local_vf_active==1) 
                   `fifo_error_check(18)                                            
              else if (local_pf_num==3 && local_vf_num=='h7ff && local_vf_active==1) 
                   `fifo_error_check(19)                                            
              else if (local_pf_num==4 && local_vf_num=='h7ff && local_vf_active==1) 
                   `fifo_error_check(20)                                           
              else if (local_pf_num==5 && local_vf_num=='h7ff && local_vf_active==1) 
                   `fifo_error_check(21)                                        
              else if (local_pf_num==6 && local_vf_num=='h7ff && local_vf_active==1) 
                   `fifo_error_check(22)                                            
              else if (local_pf_num==7 && local_vf_num=='h7ff && local_vf_active==1) 
                    `fifo_error_check(23)
              else if (local_pf_num==0 && local_vf_num==`RANDOM_VF && local_vf_active==1) 
                    `fifo_error_check(24)                                      
              else if (local_pf_num==1 && local_vf_num==`RANDOM_VF && local_vf_active==1) 
                    `fifo_error_check(25)                                      
              else if (local_pf_num==2 && local_vf_num==`RANDOM_VF && local_vf_active==1) 
                   `fifo_error_check(26)                                       
              else if (local_pf_num==3 && local_vf_num==`RANDOM_VF && local_vf_active==1) 
                   `fifo_error_check(27)                                       
              else if (local_pf_num==4 && local_vf_num==`RANDOM_VF && local_vf_active==1) 
                   `fifo_error_check(28)                                      
              else if (local_pf_num==5 && local_vf_num==`RANDOM_VF && local_vf_active==1) 
                   `fifo_error_check(29)                                   
              else if (local_pf_num==6 && local_vf_num==`RANDOM_VF && local_vf_active==1) 
                   `fifo_error_check(30)                                       
              else if (local_pf_num==7 && local_vf_num==`RANDOM_VF && local_vf_active==1) 
                    `fifo_error_check(31)

              `elsif TB_CONFIG_4
              if (local_pf_num==0 && local_vf_num==0 && local_vf_active==1) `fifo_error_check(0)
              else if (local_pf_num==0 && local_vf_num==1 && local_vf_active==1) `fifo_error_check(1)
              else if (local_pf_num==0 && local_vf_num==2 && local_vf_active==1) `fifo_error_check(2)
              else if (local_pf_num==0 && local_vf_num==3 && local_vf_active==1) `fifo_error_check(3)
              else if (local_pf_num==0 && local_vf_num==4 && local_vf_active==1) `fifo_error_check(4)
              else if (local_pf_num==0 && local_vf_num==5 && local_vf_active==1) `fifo_error_check(5)
              else if (local_pf_num==0 && local_vf_num==6 && local_vf_active==1) `fifo_error_check(6)
              else if (local_pf_num==0 && local_vf_num==7 && local_vf_active==1) `fifo_error_check(7)
              else if (local_pf_num==0 && local_vf_num==8 && local_vf_active==1) `fifo_error_check(8)
              else if (local_pf_num==0 && local_vf_num==9 && local_vf_active==1) `fifo_error_check(9)
              else if (local_pf_num==0 && local_vf_num==10 && local_vf_active==1) `fifo_error_check(10)
              else if (local_pf_num==0 && local_vf_num==11 && local_vf_active==1) `fifo_error_check(11)
              else if (local_pf_num==0 && local_vf_num==12 && local_vf_active==1) `fifo_error_check(12)
              else if (local_pf_num==0 && local_vf_num==13 && local_vf_active==1) `fifo_error_check(13)
              else if (local_pf_num==0 && local_vf_num==14 && local_vf_active==1) `fifo_error_check(14)
              else if (local_pf_num==0 && local_vf_num==15 && local_vf_active==1) `fifo_error_check(15)
              else if (local_pf_num==0 && local_vf_num==16 && local_vf_active==1) `fifo_error_check(16)
              else if (local_pf_num==0 && local_vf_num==17 && local_vf_active==1) `fifo_error_check(17)
              else if (local_pf_num==0 && local_vf_num==18 && local_vf_active==1) `fifo_error_check(18)
              else if (local_pf_num==0 && local_vf_num==19 && local_vf_active==1) `fifo_error_check(19)
              else if (local_pf_num==0 && local_vf_num==20 && local_vf_active==1) `fifo_error_check(20)
              else if (local_pf_num==0 && local_vf_num==21 && local_vf_active==1) `fifo_error_check(21)
              else if (local_pf_num==0 && local_vf_num==22 && local_vf_active==1) `fifo_error_check(22)
              else if (local_pf_num==0 && local_vf_num==23 && local_vf_active==1) `fifo_error_check(23)
              else if (local_pf_num==0 && local_vf_num==24 && local_vf_active==1) `fifo_error_check(24)
              else if (local_pf_num==0 && local_vf_num==25 && local_vf_active==1) `fifo_error_check(25)
              else if (local_pf_num==0 && local_vf_num==26 && local_vf_active==1) `fifo_error_check(26)
              else if (local_pf_num==0 && local_vf_num==27 && local_vf_active==1) `fifo_error_check(27)
              else if (local_pf_num==0 && local_vf_num==28 && local_vf_active==1) `fifo_error_check(28)
              else if (local_pf_num==0 && local_vf_num==29 && local_vf_active==1) `fifo_error_check(29)
              else if (local_pf_num==0 && local_vf_num==30 && local_vf_active==1) `fifo_error_check(30)
              else if (local_pf_num==0 && local_vf_num==31 && local_vf_active==1) `fifo_error_check(31)
              else if (local_pf_num==0 && local_vf_num==32 && local_vf_active==1) `fifo_error_check(32)
              else if (local_pf_num==0 && local_vf_num==33 && local_vf_active==1) `fifo_error_check(33)
              else if (local_pf_num==0 && local_vf_num==34 && local_vf_active==1) `fifo_error_check(34)
              else if (local_pf_num==0 && local_vf_num==35 && local_vf_active==1) `fifo_error_check(35)
              else if (local_pf_num==0 && local_vf_num==36 && local_vf_active==1) `fifo_error_check(36)
              else if (local_pf_num==0 && local_vf_num==37 && local_vf_active==1) `fifo_error_check(37)
              else if (local_pf_num==0 && local_vf_num==38 && local_vf_active==1) `fifo_error_check(38)
              else if (local_pf_num==0 && local_vf_num==39 && local_vf_active==1) `fifo_error_check(39)
              else if (local_pf_num==0 && local_vf_num==40 && local_vf_active==1) `fifo_error_check(40)
              else if (local_pf_num==0 && local_vf_num==41 && local_vf_active==1) `fifo_error_check(41)
              else if (local_pf_num==0 && local_vf_num==42 && local_vf_active==1) `fifo_error_check(42)
              else if (local_pf_num==0 && local_vf_num==43 && local_vf_active==1) `fifo_error_check(43)
              else if (local_pf_num==0 && local_vf_num==44 && local_vf_active==1) `fifo_error_check(44)
              else if (local_pf_num==0 && local_vf_num==45 && local_vf_active==1) `fifo_error_check(45)
              else if (local_pf_num==0 && local_vf_num==46 && local_vf_active==1) `fifo_error_check(46)
              else if (local_pf_num==0 && local_vf_num==47 && local_vf_active==1) `fifo_error_check(47)
              else if (local_pf_num==0 && local_vf_num==48 && local_vf_active==1) `fifo_error_check(48)
              else if (local_pf_num==0 && local_vf_num==49 && local_vf_active==1) `fifo_error_check(49)
              else if (local_pf_num==0 && local_vf_num==50 && local_vf_active==1) `fifo_error_check(50)
              else if (local_pf_num==0 && local_vf_num==51 && local_vf_active==1) `fifo_error_check(51)
              else if (local_pf_num==0 && local_vf_num==52 && local_vf_active==1) `fifo_error_check(52)
              else if (local_pf_num==0 && local_vf_num==53 && local_vf_active==1) `fifo_error_check(53)
              else if (local_pf_num==0 && local_vf_num==54 && local_vf_active==1) `fifo_error_check(54)
              else if (local_pf_num==0 && local_vf_num==55 && local_vf_active==1) `fifo_error_check(55)
              else if (local_pf_num==0 && local_vf_num==56 && local_vf_active==1) `fifo_error_check(56)
              else if (local_pf_num==0 && local_vf_num==57 && local_vf_active==1) `fifo_error_check(57)
              else if (local_pf_num==0 && local_vf_num==58 && local_vf_active==1) `fifo_error_check(58)
              else if (local_pf_num==0 && local_vf_num==59 && local_vf_active==1) `fifo_error_check(59)
              else if (local_pf_num==0 && local_vf_num==60 && local_vf_active==1) `fifo_error_check(60)
              else if (local_pf_num==0 && local_vf_num==61 && local_vf_active==1) `fifo_error_check(61)
              else if (local_pf_num==0 && local_vf_num==62 && local_vf_active==1) `fifo_error_check(62)
              else if (local_pf_num==0 && local_vf_num==63 && local_vf_active==1) `fifo_error_check(63)
              else if (local_pf_num==0 && local_vf_num==64 && local_vf_active==1) `fifo_error_check(64)
              else if (local_pf_num==0 && local_vf_num==65 && local_vf_active==1) `fifo_error_check(65)
              else if (local_pf_num==0 && local_vf_num==66 && local_vf_active==1) `fifo_error_check(66)
              else if (local_pf_num==0 && local_vf_num==67 && local_vf_active==1) `fifo_error_check(67)
              else if (local_pf_num==0 && local_vf_num==68 && local_vf_active==1) `fifo_error_check(68)
              else if (local_pf_num==0 && local_vf_num==69 && local_vf_active==1) `fifo_error_check(69)
              else if (local_pf_num==0 && local_vf_num==70 && local_vf_active==1) `fifo_error_check(70)
              else if (local_pf_num==0 && local_vf_num==71 && local_vf_active==1) `fifo_error_check(71)
              else if (local_pf_num==0 && local_vf_num==72 && local_vf_active==1) `fifo_error_check(72)
              else if (local_pf_num==0 && local_vf_num==73 && local_vf_active==1) `fifo_error_check(73)
              else if (local_pf_num==0 && local_vf_num==74 && local_vf_active==1) `fifo_error_check(74)
              else if (local_pf_num==0 && local_vf_num==75 && local_vf_active==1) `fifo_error_check(75)
              else if (local_pf_num==0 && local_vf_num==76 && local_vf_active==1) `fifo_error_check(76)
              else if (local_pf_num==0 && local_vf_num==77 && local_vf_active==1) `fifo_error_check(77)
              else if (local_pf_num==0 && local_vf_num==78 && local_vf_active==1) `fifo_error_check(78)
              else if (local_pf_num==0 && local_vf_num==79 && local_vf_active==1) `fifo_error_check(79)
              else if (local_pf_num==0 && local_vf_num==80 && local_vf_active==1) `fifo_error_check(80)
              else if (local_pf_num==0 && local_vf_num==81 && local_vf_active==1) `fifo_error_check(81)
              else if (local_pf_num==0 && local_vf_num==82 && local_vf_active==1) `fifo_error_check(82)
              else if (local_pf_num==0 && local_vf_num==83 && local_vf_active==1) `fifo_error_check(83)
              else if (local_pf_num==0 && local_vf_num==84 && local_vf_active==1) `fifo_error_check(84)
              else if (local_pf_num==0 && local_vf_num==85 && local_vf_active==1) `fifo_error_check(85)
              else if (local_pf_num==0 && local_vf_num==86 && local_vf_active==1) `fifo_error_check(86)
              else if (local_pf_num==0 && local_vf_num==87 && local_vf_active==1) `fifo_error_check(87)
              else if (local_pf_num==0 && local_vf_num==88 && local_vf_active==1) `fifo_error_check(88)
              else if (local_pf_num==0 && local_vf_num==89 && local_vf_active==1) `fifo_error_check(89)
              else if (local_pf_num==0 && local_vf_num==90 && local_vf_active==1) `fifo_error_check(90)
              else if (local_pf_num==0 && local_vf_num==91 && local_vf_active==1) `fifo_error_check(91)
              else if (local_pf_num==0 && local_vf_num==92 && local_vf_active==1) `fifo_error_check(92)
              else if (local_pf_num==0 && local_vf_num==93 && local_vf_active==1) `fifo_error_check(93)
              else if (local_pf_num==0 && local_vf_num==94 && local_vf_active==1) `fifo_error_check(94)
              else if (local_pf_num==0 && local_vf_num==95 && local_vf_active==1) `fifo_error_check(95)
              else if (local_pf_num==0 && local_vf_num==96 && local_vf_active==1) `fifo_error_check(96)
              else if (local_pf_num==0 && local_vf_num==97 && local_vf_active==1) `fifo_error_check(97)
              else if (local_pf_num==0 && local_vf_num==98 && local_vf_active==1) `fifo_error_check(98)
              else if (local_pf_num==0 && local_vf_num==99 && local_vf_active==1) `fifo_error_check(99)
              else if (local_pf_num==0 && local_vf_num==100 && local_vf_active==1) `fifo_error_check(100)
              else if (local_pf_num==0 && local_vf_num==101 && local_vf_active==1) `fifo_error_check(101)
              else if (local_pf_num==0 && local_vf_num==102 && local_vf_active==1) `fifo_error_check(102)
              else if (local_pf_num==0 && local_vf_num==103 && local_vf_active==1) `fifo_error_check(103)
              else if (local_pf_num==0 && local_vf_num==104 && local_vf_active==1) `fifo_error_check(104)
              else if (local_pf_num==0 && local_vf_num==105 && local_vf_active==1) `fifo_error_check(105)
              else if (local_pf_num==0 && local_vf_num==106 && local_vf_active==1) `fifo_error_check(106)
              else if (local_pf_num==0 && local_vf_num==107 && local_vf_active==1) `fifo_error_check(107)
              else if (local_pf_num==0 && local_vf_num==108 && local_vf_active==1) `fifo_error_check(108)
              else if (local_pf_num==0 && local_vf_num==109 && local_vf_active==1) `fifo_error_check(109)
              else if (local_pf_num==0 && local_vf_num==110 && local_vf_active==1) `fifo_error_check(110)
              else if (local_pf_num==0 && local_vf_num==111 && local_vf_active==1) `fifo_error_check(111)
              else if (local_pf_num==0 && local_vf_num==112 && local_vf_active==1) `fifo_error_check(112)
              else if (local_pf_num==0 && local_vf_num==113 && local_vf_active==1) `fifo_error_check(113)
              else if (local_pf_num==0 && local_vf_num==114 && local_vf_active==1) `fifo_error_check(114)
              else if (local_pf_num==0 && local_vf_num==115 && local_vf_active==1) `fifo_error_check(115)
              else if (local_pf_num==0 && local_vf_num==116 && local_vf_active==1) `fifo_error_check(116)
              else if (local_pf_num==0 && local_vf_num==117 && local_vf_active==1) `fifo_error_check(117)
              else if (local_pf_num==0 && local_vf_num==118 && local_vf_active==1) `fifo_error_check(118)
              else if (local_pf_num==0 && local_vf_num==119 && local_vf_active==1) `fifo_error_check(119)
              else if (local_pf_num==0 && local_vf_num==120 && local_vf_active==1) `fifo_error_check(120)
              else if (local_pf_num==0 && local_vf_num==121 && local_vf_active==1) `fifo_error_check(121)
              else if (local_pf_num==0 && local_vf_num==122 && local_vf_active==1) `fifo_error_check(122)
              else if (local_pf_num==0 && local_vf_num==123 && local_vf_active==1) `fifo_error_check(123)
              else if (local_pf_num==0 && local_vf_num==124 && local_vf_active==1) `fifo_error_check(124)
              else if (local_pf_num==0 && local_vf_num==125 && local_vf_active==1) `fifo_error_check(125)
              else if (local_pf_num==0 && local_vf_num==126 && local_vf_active==1) `fifo_error_check(126)
              else if (local_pf_num==0 && local_vf_num==127 && local_vf_active==1) `fifo_error_check(127)
              else if (local_pf_num==0 && local_vf_num==128 && local_vf_active==1) `fifo_error_check(128)
              else if (local_pf_num==0 && local_vf_num==129 && local_vf_active==1) `fifo_error_check(129)
              else if (local_pf_num==0 && local_vf_num==130 && local_vf_active==1) `fifo_error_check(130)
              else if (local_pf_num==0 && local_vf_num==131 && local_vf_active==1) `fifo_error_check(131)
              else if (local_pf_num==0 && local_vf_num==132 && local_vf_active==1) `fifo_error_check(132)
              else if (local_pf_num==0 && local_vf_num==133 && local_vf_active==1) `fifo_error_check(133)
              else if (local_pf_num==0 && local_vf_num==134 && local_vf_active==1) `fifo_error_check(134)
              else if (local_pf_num==0 && local_vf_num==135 && local_vf_active==1) `fifo_error_check(135)
              else if (local_pf_num==0 && local_vf_num==136 && local_vf_active==1) `fifo_error_check(136)
              else if (local_pf_num==0 && local_vf_num==137 && local_vf_active==1) `fifo_error_check(137)
              else if (local_pf_num==0 && local_vf_num==138 && local_vf_active==1) `fifo_error_check(138)
              else if (local_pf_num==0 && local_vf_num==139 && local_vf_active==1) `fifo_error_check(139)
              else if (local_pf_num==0 && local_vf_num==140 && local_vf_active==1) `fifo_error_check(140)
              else if (local_pf_num==0 && local_vf_num==141 && local_vf_active==1) `fifo_error_check(141)
              else if (local_pf_num==0 && local_vf_num==142 && local_vf_active==1) `fifo_error_check(142)
              else if (local_pf_num==0 && local_vf_num==143 && local_vf_active==1) `fifo_error_check(143)
              else if (local_pf_num==0 && local_vf_num==144 && local_vf_active==1) `fifo_error_check(144)
              else if (local_pf_num==0 && local_vf_num==145 && local_vf_active==1) `fifo_error_check(145)
              else if (local_pf_num==0 && local_vf_num==146 && local_vf_active==1) `fifo_error_check(146)
              else if (local_pf_num==0 && local_vf_num==147 && local_vf_active==1) `fifo_error_check(147)
              else if (local_pf_num==0 && local_vf_num==148 && local_vf_active==1) `fifo_error_check(148)
              else if (local_pf_num==0 && local_vf_num==149 && local_vf_active==1) `fifo_error_check(149)
              else if (local_pf_num==0 && local_vf_num==150 && local_vf_active==1) `fifo_error_check(150)
              else if (local_pf_num==0 && local_vf_num==151 && local_vf_active==1) `fifo_error_check(151)
              else if (local_pf_num==0 && local_vf_num==152 && local_vf_active==1) `fifo_error_check(152)
              else if (local_pf_num==0 && local_vf_num==153 && local_vf_active==1) `fifo_error_check(153)
              else if (local_pf_num==0 && local_vf_num==154 && local_vf_active==1) `fifo_error_check(154)
              else if (local_pf_num==0 && local_vf_num==155 && local_vf_active==1) `fifo_error_check(155)
              else if (local_pf_num==0 && local_vf_num==156 && local_vf_active==1) `fifo_error_check(156)
              else if (local_pf_num==0 && local_vf_num==157 && local_vf_active==1) `fifo_error_check(157)
              else if (local_pf_num==0 && local_vf_num==158 && local_vf_active==1) `fifo_error_check(158)
              else if (local_pf_num==0 && local_vf_num==159 && local_vf_active==1) `fifo_error_check(159)
              else if (local_pf_num==0 && local_vf_num==160 && local_vf_active==1) `fifo_error_check(160)
              else if (local_pf_num==0 && local_vf_num==161 && local_vf_active==1) `fifo_error_check(161)
              else if (local_pf_num==0 && local_vf_num==162 && local_vf_active==1) `fifo_error_check(162)
              else if (local_pf_num==0 && local_vf_num==163 && local_vf_active==1) `fifo_error_check(163)
              else if (local_pf_num==0 && local_vf_num==164 && local_vf_active==1) `fifo_error_check(164)
              else if (local_pf_num==0 && local_vf_num==165 && local_vf_active==1) `fifo_error_check(165)
              else if (local_pf_num==0 && local_vf_num==166 && local_vf_active==1) `fifo_error_check(166)
              else if (local_pf_num==0 && local_vf_num==167 && local_vf_active==1) `fifo_error_check(167)
              else if (local_pf_num==0 && local_vf_num==168 && local_vf_active==1) `fifo_error_check(168)
              else if (local_pf_num==0 && local_vf_num==169 && local_vf_active==1) `fifo_error_check(169)
              else if (local_pf_num==0 && local_vf_num==170 && local_vf_active==1) `fifo_error_check(170)
              else if (local_pf_num==0 && local_vf_num==171 && local_vf_active==1) `fifo_error_check(171)
              else if (local_pf_num==0 && local_vf_num==172 && local_vf_active==1) `fifo_error_check(172)
              else if (local_pf_num==0 && local_vf_num==173 && local_vf_active==1) `fifo_error_check(173)
              else if (local_pf_num==0 && local_vf_num==174 && local_vf_active==1) `fifo_error_check(174)
              else if (local_pf_num==0 && local_vf_num==175 && local_vf_active==1) `fifo_error_check(175)
              else if (local_pf_num==0 && local_vf_num==176 && local_vf_active==1) `fifo_error_check(176)
              else if (local_pf_num==0 && local_vf_num==177 && local_vf_active==1) `fifo_error_check(177)
              else if (local_pf_num==0 && local_vf_num==178 && local_vf_active==1) `fifo_error_check(178)
              else if (local_pf_num==0 && local_vf_num==179 && local_vf_active==1) `fifo_error_check(179)
              else if (local_pf_num==0 && local_vf_num==180 && local_vf_active==1) `fifo_error_check(180)
              else if (local_pf_num==0 && local_vf_num==181 && local_vf_active==1) `fifo_error_check(181)
              else if (local_pf_num==0 && local_vf_num==182 && local_vf_active==1) `fifo_error_check(182)
              else if (local_pf_num==0 && local_vf_num==183 && local_vf_active==1) `fifo_error_check(183)
              else if (local_pf_num==0 && local_vf_num==184 && local_vf_active==1) `fifo_error_check(184)
              else if (local_pf_num==0 && local_vf_num==185 && local_vf_active==1) `fifo_error_check(185)
              else if (local_pf_num==0 && local_vf_num==186 && local_vf_active==1) `fifo_error_check(186)
              else if (local_pf_num==0 && local_vf_num==187 && local_vf_active==1) `fifo_error_check(187)
              else if (local_pf_num==0 && local_vf_num==188 && local_vf_active==1) `fifo_error_check(188)
              else if (local_pf_num==0 && local_vf_num==189 && local_vf_active==1) `fifo_error_check(189)
              else if (local_pf_num==0 && local_vf_num==190 && local_vf_active==1) `fifo_error_check(190)
              else if (local_pf_num==0 && local_vf_num==191 && local_vf_active==1) `fifo_error_check(191)
              else if (local_pf_num==0 && local_vf_num==192 && local_vf_active==1) `fifo_error_check(192)
              else if (local_pf_num==0 && local_vf_num==193 && local_vf_active==1) `fifo_error_check(193)
              else if (local_pf_num==0 && local_vf_num==194 && local_vf_active==1) `fifo_error_check(194)
              else if (local_pf_num==0 && local_vf_num==195 && local_vf_active==1) `fifo_error_check(195)
              else if (local_pf_num==0 && local_vf_num==196 && local_vf_active==1) `fifo_error_check(196)
              else if (local_pf_num==0 && local_vf_num==197 && local_vf_active==1) `fifo_error_check(197)
              else if (local_pf_num==0 && local_vf_num==198 && local_vf_active==1) `fifo_error_check(198)
              else if (local_pf_num==0 && local_vf_num==199 && local_vf_active==1) `fifo_error_check(199)
              else if (local_pf_num==0 && local_vf_num==200 && local_vf_active==1) `fifo_error_check(200)
              else if (local_pf_num==0 && local_vf_num==201 && local_vf_active==1) `fifo_error_check(201)
              else if (local_pf_num==0 && local_vf_num==202 && local_vf_active==1) `fifo_error_check(202)
              else if (local_pf_num==0 && local_vf_num==203 && local_vf_active==1) `fifo_error_check(203)
              else if (local_pf_num==0 && local_vf_num==204 && local_vf_active==1) `fifo_error_check(204)
              else if (local_pf_num==0 && local_vf_num==205 && local_vf_active==1) `fifo_error_check(205)
              else if (local_pf_num==0 && local_vf_num==206 && local_vf_active==1) `fifo_error_check(206)
              else if (local_pf_num==0 && local_vf_num==207 && local_vf_active==1) `fifo_error_check(207)
              else if (local_pf_num==0 && local_vf_num==208 && local_vf_active==1) `fifo_error_check(208)
              else if (local_pf_num==0 && local_vf_num==209 && local_vf_active==1) `fifo_error_check(209)
              else if (local_pf_num==0 && local_vf_num==210 && local_vf_active==1) `fifo_error_check(210)
              else if (local_pf_num==0 && local_vf_num==211 && local_vf_active==1) `fifo_error_check(211)
              else if (local_pf_num==0 && local_vf_num==212 && local_vf_active==1) `fifo_error_check(212)
              else if (local_pf_num==0 && local_vf_num==213 && local_vf_active==1) `fifo_error_check(213)
              else if (local_pf_num==0 && local_vf_num==214 && local_vf_active==1) `fifo_error_check(214)
              else if (local_pf_num==0 && local_vf_num==215 && local_vf_active==1) `fifo_error_check(215)
              else if (local_pf_num==0 && local_vf_num==216 && local_vf_active==1) `fifo_error_check(216)
              else if (local_pf_num==0 && local_vf_num==217 && local_vf_active==1) `fifo_error_check(217)
              else if (local_pf_num==0 && local_vf_num==218 && local_vf_active==1) `fifo_error_check(218)
              else if (local_pf_num==0 && local_vf_num==219 && local_vf_active==1) `fifo_error_check(219)
              else if (local_pf_num==0 && local_vf_num==220 && local_vf_active==1) `fifo_error_check(220)
              else if (local_pf_num==0 && local_vf_num==221 && local_vf_active==1) `fifo_error_check(221)
              else if (local_pf_num==0 && local_vf_num==222 && local_vf_active==1) `fifo_error_check(222)
              else if (local_pf_num==0 && local_vf_num==223 && local_vf_active==1) `fifo_error_check(223)
              else if (local_pf_num==0 && local_vf_num==224 && local_vf_active==1) `fifo_error_check(224)
              else if (local_pf_num==0 && local_vf_num==225 && local_vf_active==1) `fifo_error_check(225)
              else if (local_pf_num==0 && local_vf_num==226 && local_vf_active==1) `fifo_error_check(226)
              else if (local_pf_num==0 && local_vf_num==227 && local_vf_active==1) `fifo_error_check(227)
              else if (local_pf_num==0 && local_vf_num==228 && local_vf_active==1) `fifo_error_check(228)
              else if (local_pf_num==0 && local_vf_num==229 && local_vf_active==1) `fifo_error_check(229)
              else if (local_pf_num==0 && local_vf_num==230 && local_vf_active==1) `fifo_error_check(230)
              else if (local_pf_num==0 && local_vf_num==231 && local_vf_active==1) `fifo_error_check(231)
              else if (local_pf_num==0 && local_vf_num==232 && local_vf_active==1) `fifo_error_check(232)
              else if (local_pf_num==0 && local_vf_num==233 && local_vf_active==1) `fifo_error_check(233)
              else if (local_pf_num==0 && local_vf_num==234 && local_vf_active==1) `fifo_error_check(234)
              else if (local_pf_num==0 && local_vf_num==235 && local_vf_active==1) `fifo_error_check(235)
              else if (local_pf_num==0 && local_vf_num==236 && local_vf_active==1) `fifo_error_check(236)
              else if (local_pf_num==0 && local_vf_num==237 && local_vf_active==1) `fifo_error_check(237)
              else if (local_pf_num==0 && local_vf_num==238 && local_vf_active==1) `fifo_error_check(238)
              else if (local_pf_num==0 && local_vf_num==239 && local_vf_active==1) `fifo_error_check(239)
              else if (local_pf_num==0 && local_vf_num==240 && local_vf_active==1) `fifo_error_check(240)
              else if (local_pf_num==0 && local_vf_num==241 && local_vf_active==1) `fifo_error_check(241)
              else if (local_pf_num==0 && local_vf_num==242 && local_vf_active==1) `fifo_error_check(242)
              else if (local_pf_num==0 && local_vf_num==243 && local_vf_active==1) `fifo_error_check(243)
              else if (local_pf_num==0 && local_vf_num==244 && local_vf_active==1) `fifo_error_check(244)
              else if (local_pf_num==0 && local_vf_num==245 && local_vf_active==1) `fifo_error_check(245)
              else if (local_pf_num==0 && local_vf_num==246 && local_vf_active==1) `fifo_error_check(246)
              else if (local_pf_num==0 && local_vf_num==247 && local_vf_active==1) `fifo_error_check(247)
              else if (local_pf_num==0 && local_vf_num==248 && local_vf_active==1) `fifo_error_check(248)
              else if (local_pf_num==0 && local_vf_num==249 && local_vf_active==1) `fifo_error_check(249)
              else if (local_pf_num==0 && local_vf_num==250 && local_vf_active==1) `fifo_error_check(250)
              else if (local_pf_num==0 && local_vf_num==251 && local_vf_active==1) `fifo_error_check(251)
              else if (local_pf_num==0 && local_vf_num==252 && local_vf_active==1) `fifo_error_check(252)
              else if (local_pf_num==0 && local_vf_num==253 && local_vf_active==1) `fifo_error_check(253)
              else if (local_pf_num==0 && local_vf_num==254 && local_vf_active==1) `fifo_error_check(254)
              else if (local_pf_num==0 && local_vf_num==255 && local_vf_active==1) `fifo_error_check(255)
              else if (local_pf_num==0 && local_vf_num==256 && local_vf_active==1) `fifo_error_check(256)
              else if (local_pf_num==0 && local_vf_num==257 && local_vf_active==1) `fifo_error_check(257)
              else if (local_pf_num==0 && local_vf_num==258 && local_vf_active==1) `fifo_error_check(258)
              else if (local_pf_num==0 && local_vf_num==259 && local_vf_active==1) `fifo_error_check(259)
              else if (local_pf_num==0 && local_vf_num==260 && local_vf_active==1) `fifo_error_check(260)
              else if (local_pf_num==0 && local_vf_num==261 && local_vf_active==1) `fifo_error_check(261)
              else if (local_pf_num==0 && local_vf_num==262 && local_vf_active==1) `fifo_error_check(262)
              else if (local_pf_num==0 && local_vf_num==263 && local_vf_active==1) `fifo_error_check(263)
              else if (local_pf_num==0 && local_vf_num==264 && local_vf_active==1) `fifo_error_check(264)
              else if (local_pf_num==0 && local_vf_num==265 && local_vf_active==1) `fifo_error_check(265)
              else if (local_pf_num==0 && local_vf_num==266 && local_vf_active==1) `fifo_error_check(266)
              else if (local_pf_num==0 && local_vf_num==267 && local_vf_active==1) `fifo_error_check(267)
              else if (local_pf_num==0 && local_vf_num==268 && local_vf_active==1) `fifo_error_check(268)
              else if (local_pf_num==0 && local_vf_num==269 && local_vf_active==1) `fifo_error_check(269)
              else if (local_pf_num==0 && local_vf_num==270 && local_vf_active==1) `fifo_error_check(270)
              else if (local_pf_num==0 && local_vf_num==271 && local_vf_active==1) `fifo_error_check(271)
              else if (local_pf_num==0 && local_vf_num==272 && local_vf_active==1) `fifo_error_check(272)
              else if (local_pf_num==0 && local_vf_num==273 && local_vf_active==1) `fifo_error_check(273)
              else if (local_pf_num==0 && local_vf_num==274 && local_vf_active==1) `fifo_error_check(274)
              else if (local_pf_num==0 && local_vf_num==275 && local_vf_active==1) `fifo_error_check(275)
              else if (local_pf_num==0 && local_vf_num==276 && local_vf_active==1) `fifo_error_check(276)
              else if (local_pf_num==0 && local_vf_num==277 && local_vf_active==1) `fifo_error_check(277)
              else if (local_pf_num==0 && local_vf_num==278 && local_vf_active==1) `fifo_error_check(278)
              else if (local_pf_num==0 && local_vf_num==279 && local_vf_active==1) `fifo_error_check(279)
              else if (local_pf_num==0 && local_vf_num==280 && local_vf_active==1) `fifo_error_check(280)
              else if (local_pf_num==0 && local_vf_num==281 && local_vf_active==1) `fifo_error_check(281)
              else if (local_pf_num==0 && local_vf_num==282 && local_vf_active==1) `fifo_error_check(282)
              else if (local_pf_num==0 && local_vf_num==283 && local_vf_active==1) `fifo_error_check(283)
              else if (local_pf_num==0 && local_vf_num==284 && local_vf_active==1) `fifo_error_check(284)
              else if (local_pf_num==0 && local_vf_num==285 && local_vf_active==1) `fifo_error_check(285)
              else if (local_pf_num==0 && local_vf_num==286 && local_vf_active==1) `fifo_error_check(286)
              else if (local_pf_num==0 && local_vf_num==287 && local_vf_active==1) `fifo_error_check(287)
              else if (local_pf_num==0 && local_vf_num==288 && local_vf_active==1) `fifo_error_check(288)
              else if (local_pf_num==0 && local_vf_num==289 && local_vf_active==1) `fifo_error_check(289)
              else if (local_pf_num==0 && local_vf_num==290 && local_vf_active==1) `fifo_error_check(290)
              else if (local_pf_num==0 && local_vf_num==291 && local_vf_active==1) `fifo_error_check(291)
              else if (local_pf_num==0 && local_vf_num==292 && local_vf_active==1) `fifo_error_check(292)
              else if (local_pf_num==0 && local_vf_num==293 && local_vf_active==1) `fifo_error_check(293)
              else if (local_pf_num==0 && local_vf_num==294 && local_vf_active==1) `fifo_error_check(294)
              else if (local_pf_num==0 && local_vf_num==295 && local_vf_active==1) `fifo_error_check(295)
              else if (local_pf_num==0 && local_vf_num==296 && local_vf_active==1) `fifo_error_check(296)
              else if (local_pf_num==0 && local_vf_num==297 && local_vf_active==1) `fifo_error_check(297)
              else if (local_pf_num==0 && local_vf_num==298 && local_vf_active==1) `fifo_error_check(298)
              else if (local_pf_num==0 && local_vf_num==299 && local_vf_active==1) `fifo_error_check(299)
              else if (local_pf_num==0 && local_vf_num==300 && local_vf_active==1) `fifo_error_check(300)
              else if (local_pf_num==0 && local_vf_num==301 && local_vf_active==1) `fifo_error_check(301)
              else if (local_pf_num==0 && local_vf_num==302 && local_vf_active==1) `fifo_error_check(302)
              else if (local_pf_num==0 && local_vf_num==303 && local_vf_active==1) `fifo_error_check(303)
              else if (local_pf_num==0 && local_vf_num==304 && local_vf_active==1) `fifo_error_check(304)
              else if (local_pf_num==0 && local_vf_num==305 && local_vf_active==1) `fifo_error_check(305)
              else if (local_pf_num==0 && local_vf_num==306 && local_vf_active==1) `fifo_error_check(306)
              else if (local_pf_num==0 && local_vf_num==307 && local_vf_active==1) `fifo_error_check(307)
              else if (local_pf_num==0 && local_vf_num==308 && local_vf_active==1) `fifo_error_check(308)
              else if (local_pf_num==0 && local_vf_num==309 && local_vf_active==1) `fifo_error_check(309)
              else if (local_pf_num==0 && local_vf_num==310 && local_vf_active==1) `fifo_error_check(310)
              else if (local_pf_num==0 && local_vf_num==311 && local_vf_active==1) `fifo_error_check(311)
              else if (local_pf_num==0 && local_vf_num==312 && local_vf_active==1) `fifo_error_check(312)
              else if (local_pf_num==0 && local_vf_num==313 && local_vf_active==1) `fifo_error_check(313)
              else if (local_pf_num==0 && local_vf_num==314 && local_vf_active==1) `fifo_error_check(314)
              else if (local_pf_num==0 && local_vf_num==315 && local_vf_active==1) `fifo_error_check(315)
              else if (local_pf_num==0 && local_vf_num==316 && local_vf_active==1) `fifo_error_check(316)
              else if (local_pf_num==0 && local_vf_num==317 && local_vf_active==1) `fifo_error_check(317)
              else if (local_pf_num==0 && local_vf_num==318 && local_vf_active==1) `fifo_error_check(318)
              else if (local_pf_num==0 && local_vf_num==319 && local_vf_active==1) `fifo_error_check(319)
              else if (local_pf_num==0 && local_vf_num==320 && local_vf_active==1) `fifo_error_check(320)
              else if (local_pf_num==0 && local_vf_num==321 && local_vf_active==1) `fifo_error_check(321)
              else if (local_pf_num==0 && local_vf_num==322 && local_vf_active==1) `fifo_error_check(322)
              else if (local_pf_num==0 && local_vf_num==323 && local_vf_active==1) `fifo_error_check(323)
              else if (local_pf_num==0 && local_vf_num==324 && local_vf_active==1) `fifo_error_check(324)
              else if (local_pf_num==0 && local_vf_num==325 && local_vf_active==1) `fifo_error_check(325)
              else if (local_pf_num==0 && local_vf_num==326 && local_vf_active==1) `fifo_error_check(326)
              else if (local_pf_num==0 && local_vf_num==327 && local_vf_active==1) `fifo_error_check(327)
              else if (local_pf_num==0 && local_vf_num==328 && local_vf_active==1) `fifo_error_check(328)
              else if (local_pf_num==0 && local_vf_num==329 && local_vf_active==1) `fifo_error_check(329)
              else if (local_pf_num==0 && local_vf_num==330 && local_vf_active==1) `fifo_error_check(330)
              else if (local_pf_num==0 && local_vf_num==331 && local_vf_active==1) `fifo_error_check(331)
              else if (local_pf_num==0 && local_vf_num==332 && local_vf_active==1) `fifo_error_check(332)
              else if (local_pf_num==0 && local_vf_num==333 && local_vf_active==1) `fifo_error_check(333)
              else if (local_pf_num==0 && local_vf_num==334 && local_vf_active==1) `fifo_error_check(334)
              else if (local_pf_num==0 && local_vf_num==335 && local_vf_active==1) `fifo_error_check(335)
              else if (local_pf_num==0 && local_vf_num==336 && local_vf_active==1) `fifo_error_check(336)
              else if (local_pf_num==0 && local_vf_num==337 && local_vf_active==1) `fifo_error_check(337)
              else if (local_pf_num==0 && local_vf_num==338 && local_vf_active==1) `fifo_error_check(338)
              else if (local_pf_num==0 && local_vf_num==339 && local_vf_active==1) `fifo_error_check(339)
              else if (local_pf_num==0 && local_vf_num==340 && local_vf_active==1) `fifo_error_check(340)
              else if (local_pf_num==0 && local_vf_num==341 && local_vf_active==1) `fifo_error_check(341)
              else if (local_pf_num==0 && local_vf_num==342 && local_vf_active==1) `fifo_error_check(342)
              else if (local_pf_num==0 && local_vf_num==343 && local_vf_active==1) `fifo_error_check(343)
              else if (local_pf_num==0 && local_vf_num==344 && local_vf_active==1) `fifo_error_check(344)
              else if (local_pf_num==0 && local_vf_num==345 && local_vf_active==1) `fifo_error_check(345)
              else if (local_pf_num==0 && local_vf_num==346 && local_vf_active==1) `fifo_error_check(346)
              else if (local_pf_num==0 && local_vf_num==347 && local_vf_active==1) `fifo_error_check(347)
              else if (local_pf_num==0 && local_vf_num==348 && local_vf_active==1) `fifo_error_check(348)
              else if (local_pf_num==0 && local_vf_num==349 && local_vf_active==1) `fifo_error_check(349)
              else if (local_pf_num==0 && local_vf_num==350 && local_vf_active==1) `fifo_error_check(350)
              else if (local_pf_num==0 && local_vf_num==351 && local_vf_active==1) `fifo_error_check(351)
              else if (local_pf_num==0 && local_vf_num==352 && local_vf_active==1) `fifo_error_check(352)
              else if (local_pf_num==0 && local_vf_num==353 && local_vf_active==1) `fifo_error_check(353)
              else if (local_pf_num==0 && local_vf_num==354 && local_vf_active==1) `fifo_error_check(354)
              else if (local_pf_num==0 && local_vf_num==355 && local_vf_active==1) `fifo_error_check(355)
              else if (local_pf_num==0 && local_vf_num==356 && local_vf_active==1) `fifo_error_check(356)
              else if (local_pf_num==0 && local_vf_num==357 && local_vf_active==1) `fifo_error_check(357)
              else if (local_pf_num==0 && local_vf_num==358 && local_vf_active==1) `fifo_error_check(358)
              else if (local_pf_num==0 && local_vf_num==359 && local_vf_active==1) `fifo_error_check(359)
              else if (local_pf_num==0 && local_vf_num==360 && local_vf_active==1) `fifo_error_check(360)
              else if (local_pf_num==0 && local_vf_num==361 && local_vf_active==1) `fifo_error_check(361)
              else if (local_pf_num==0 && local_vf_num==362 && local_vf_active==1) `fifo_error_check(362)
              else if (local_pf_num==0 && local_vf_num==363 && local_vf_active==1) `fifo_error_check(363)
              else if (local_pf_num==0 && local_vf_num==364 && local_vf_active==1) `fifo_error_check(364)
              else if (local_pf_num==0 && local_vf_num==365 && local_vf_active==1) `fifo_error_check(365)
              else if (local_pf_num==0 && local_vf_num==366 && local_vf_active==1) `fifo_error_check(366)
              else if (local_pf_num==0 && local_vf_num==367 && local_vf_active==1) `fifo_error_check(367)
              else if (local_pf_num==0 && local_vf_num==368 && local_vf_active==1) `fifo_error_check(368)
              else if (local_pf_num==0 && local_vf_num==369 && local_vf_active==1) `fifo_error_check(369)
              else if (local_pf_num==0 && local_vf_num==370 && local_vf_active==1) `fifo_error_check(370)
              else if (local_pf_num==0 && local_vf_num==371 && local_vf_active==1) `fifo_error_check(371)
              else if (local_pf_num==0 && local_vf_num==372 && local_vf_active==1) `fifo_error_check(372)
              else if (local_pf_num==0 && local_vf_num==373 && local_vf_active==1) `fifo_error_check(373)
              else if (local_pf_num==0 && local_vf_num==374 && local_vf_active==1) `fifo_error_check(374)
              else if (local_pf_num==0 && local_vf_num==375 && local_vf_active==1) `fifo_error_check(375)
              else if (local_pf_num==0 && local_vf_num==376 && local_vf_active==1) `fifo_error_check(376)
              else if (local_pf_num==0 && local_vf_num==377 && local_vf_active==1) `fifo_error_check(377)
              else if (local_pf_num==0 && local_vf_num==378 && local_vf_active==1) `fifo_error_check(378)
              else if (local_pf_num==0 && local_vf_num==379 && local_vf_active==1) `fifo_error_check(379)
              else if (local_pf_num==0 && local_vf_num==380 && local_vf_active==1) `fifo_error_check(380)
              else if (local_pf_num==0 && local_vf_num==381 && local_vf_active==1) `fifo_error_check(381)
              else if (local_pf_num==0 && local_vf_num==382 && local_vf_active==1) `fifo_error_check(382)
              else if (local_pf_num==0 && local_vf_num==383 && local_vf_active==1) `fifo_error_check(383)
              else if (local_pf_num==0 && local_vf_num==384 && local_vf_active==1) `fifo_error_check(384)
              else if (local_pf_num==0 && local_vf_num==385 && local_vf_active==1) `fifo_error_check(385)
              else if (local_pf_num==0 && local_vf_num==386 && local_vf_active==1) `fifo_error_check(386)
              else if (local_pf_num==0 && local_vf_num==387 && local_vf_active==1) `fifo_error_check(387)
              else if (local_pf_num==0 && local_vf_num==388 && local_vf_active==1) `fifo_error_check(388)
              else if (local_pf_num==0 && local_vf_num==389 && local_vf_active==1) `fifo_error_check(389)
              else if (local_pf_num==0 && local_vf_num==390 && local_vf_active==1) `fifo_error_check(390)
              else if (local_pf_num==0 && local_vf_num==391 && local_vf_active==1) `fifo_error_check(391)
              else if (local_pf_num==0 && local_vf_num==392 && local_vf_active==1) `fifo_error_check(392)
              else if (local_pf_num==0 && local_vf_num==393 && local_vf_active==1) `fifo_error_check(393)
              else if (local_pf_num==0 && local_vf_num==394 && local_vf_active==1) `fifo_error_check(394)
              else if (local_pf_num==0 && local_vf_num==395 && local_vf_active==1) `fifo_error_check(395)
              else if (local_pf_num==0 && local_vf_num==396 && local_vf_active==1) `fifo_error_check(396)
              else if (local_pf_num==0 && local_vf_num==397 && local_vf_active==1) `fifo_error_check(397)
              else if (local_pf_num==0 && local_vf_num==398 && local_vf_active==1) `fifo_error_check(398)
              else if (local_pf_num==0 && local_vf_num==399 && local_vf_active==1) `fifo_error_check(399)
              else if (local_pf_num==0 && local_vf_num==400 && local_vf_active==1) `fifo_error_check(400)
              else if (local_pf_num==0 && local_vf_num==401 && local_vf_active==1) `fifo_error_check(401)
              else if (local_pf_num==0 && local_vf_num==402 && local_vf_active==1) `fifo_error_check(402)
              else if (local_pf_num==0 && local_vf_num==403 && local_vf_active==1) `fifo_error_check(403)
              else if (local_pf_num==0 && local_vf_num==404 && local_vf_active==1) `fifo_error_check(404)
              else if (local_pf_num==0 && local_vf_num==405 && local_vf_active==1) `fifo_error_check(405)
              else if (local_pf_num==0 && local_vf_num==406 && local_vf_active==1) `fifo_error_check(406)
              else if (local_pf_num==0 && local_vf_num==407 && local_vf_active==1) `fifo_error_check(407)
              else if (local_pf_num==0 && local_vf_num==408 && local_vf_active==1) `fifo_error_check(408)
              else if (local_pf_num==0 && local_vf_num==409 && local_vf_active==1) `fifo_error_check(409)
              else if (local_pf_num==0 && local_vf_num==410 && local_vf_active==1) `fifo_error_check(410)
              else if (local_pf_num==0 && local_vf_num==411 && local_vf_active==1) `fifo_error_check(411)
              else if (local_pf_num==0 && local_vf_num==412 && local_vf_active==1) `fifo_error_check(412)
              else if (local_pf_num==0 && local_vf_num==413 && local_vf_active==1) `fifo_error_check(413)
              else if (local_pf_num==0 && local_vf_num==414 && local_vf_active==1) `fifo_error_check(414)
              else if (local_pf_num==0 && local_vf_num==415 && local_vf_active==1) `fifo_error_check(415)
              else if (local_pf_num==0 && local_vf_num==416 && local_vf_active==1) `fifo_error_check(416)
              else if (local_pf_num==0 && local_vf_num==417 && local_vf_active==1) `fifo_error_check(417)
              else if (local_pf_num==0 && local_vf_num==418 && local_vf_active==1) `fifo_error_check(418)
              else if (local_pf_num==0 && local_vf_num==419 && local_vf_active==1) `fifo_error_check(419)
              else if (local_pf_num==0 && local_vf_num==420 && local_vf_active==1) `fifo_error_check(420)
              else if (local_pf_num==0 && local_vf_num==421 && local_vf_active==1) `fifo_error_check(421)
              else if (local_pf_num==0 && local_vf_num==422 && local_vf_active==1) `fifo_error_check(422)
              else if (local_pf_num==0 && local_vf_num==423 && local_vf_active==1) `fifo_error_check(423)
              else if (local_pf_num==0 && local_vf_num==424 && local_vf_active==1) `fifo_error_check(424)
              else if (local_pf_num==0 && local_vf_num==425 && local_vf_active==1) `fifo_error_check(425)
              else if (local_pf_num==0 && local_vf_num==426 && local_vf_active==1) `fifo_error_check(426)
              else if (local_pf_num==0 && local_vf_num==427 && local_vf_active==1) `fifo_error_check(427)
              else if (local_pf_num==0 && local_vf_num==428 && local_vf_active==1) `fifo_error_check(428)
              else if (local_pf_num==0 && local_vf_num==429 && local_vf_active==1) `fifo_error_check(429)
              else if (local_pf_num==0 && local_vf_num==430 && local_vf_active==1) `fifo_error_check(430)
              else if (local_pf_num==0 && local_vf_num==431 && local_vf_active==1) `fifo_error_check(431)
              else if (local_pf_num==0 && local_vf_num==432 && local_vf_active==1) `fifo_error_check(432)
              else if (local_pf_num==0 && local_vf_num==433 && local_vf_active==1) `fifo_error_check(433)
              else if (local_pf_num==0 && local_vf_num==434 && local_vf_active==1) `fifo_error_check(434)
              else if (local_pf_num==0 && local_vf_num==435 && local_vf_active==1) `fifo_error_check(435)
              else if (local_pf_num==0 && local_vf_num==436 && local_vf_active==1) `fifo_error_check(436)
              else if (local_pf_num==0 && local_vf_num==437 && local_vf_active==1) `fifo_error_check(437)
              else if (local_pf_num==0 && local_vf_num==438 && local_vf_active==1) `fifo_error_check(438)
              else if (local_pf_num==0 && local_vf_num==439 && local_vf_active==1) `fifo_error_check(439)
              else if (local_pf_num==0 && local_vf_num==440 && local_vf_active==1) `fifo_error_check(440)
              else if (local_pf_num==0 && local_vf_num==441 && local_vf_active==1) `fifo_error_check(441)
              else if (local_pf_num==0 && local_vf_num==442 && local_vf_active==1) `fifo_error_check(442)
              else if (local_pf_num==0 && local_vf_num==443 && local_vf_active==1) `fifo_error_check(443)
              else if (local_pf_num==0 && local_vf_num==444 && local_vf_active==1) `fifo_error_check(444)
              else if (local_pf_num==0 && local_vf_num==445 && local_vf_active==1) `fifo_error_check(445)
              else if (local_pf_num==0 && local_vf_num==446 && local_vf_active==1) `fifo_error_check(446)
              else if (local_pf_num==0 && local_vf_num==447 && local_vf_active==1) `fifo_error_check(447)
              else if (local_pf_num==0 && local_vf_num==448 && local_vf_active==1) `fifo_error_check(448)
              else if (local_pf_num==0 && local_vf_num==449 && local_vf_active==1) `fifo_error_check(449)
              else if (local_pf_num==0 && local_vf_num==450 && local_vf_active==1) `fifo_error_check(450)
              else if (local_pf_num==0 && local_vf_num==451 && local_vf_active==1) `fifo_error_check(451)
              else if (local_pf_num==0 && local_vf_num==452 && local_vf_active==1) `fifo_error_check(452)
              else if (local_pf_num==0 && local_vf_num==453 && local_vf_active==1) `fifo_error_check(453)
              else if (local_pf_num==0 && local_vf_num==454 && local_vf_active==1) `fifo_error_check(454)
              else if (local_pf_num==0 && local_vf_num==455 && local_vf_active==1) `fifo_error_check(455)
              else if (local_pf_num==0 && local_vf_num==456 && local_vf_active==1) `fifo_error_check(456)
              else if (local_pf_num==0 && local_vf_num==457 && local_vf_active==1) `fifo_error_check(457)
              else if (local_pf_num==0 && local_vf_num==458 && local_vf_active==1) `fifo_error_check(458)
              else if (local_pf_num==0 && local_vf_num==459 && local_vf_active==1) `fifo_error_check(459)
              else if (local_pf_num==0 && local_vf_num==460 && local_vf_active==1) `fifo_error_check(460)
              else if (local_pf_num==0 && local_vf_num==461 && local_vf_active==1) `fifo_error_check(461)
              else if (local_pf_num==0 && local_vf_num==462 && local_vf_active==1) `fifo_error_check(462)
              else if (local_pf_num==0 && local_vf_num==463 && local_vf_active==1) `fifo_error_check(463)
              else if (local_pf_num==0 && local_vf_num==464 && local_vf_active==1) `fifo_error_check(464)
              else if (local_pf_num==0 && local_vf_num==465 && local_vf_active==1) `fifo_error_check(465)
              else if (local_pf_num==0 && local_vf_num==466 && local_vf_active==1) `fifo_error_check(466)
              else if (local_pf_num==0 && local_vf_num==467 && local_vf_active==1) `fifo_error_check(467)
              else if (local_pf_num==0 && local_vf_num==468 && local_vf_active==1) `fifo_error_check(468)
              else if (local_pf_num==0 && local_vf_num==469 && local_vf_active==1) `fifo_error_check(469)
              else if (local_pf_num==0 && local_vf_num==470 && local_vf_active==1) `fifo_error_check(470)
              else if (local_pf_num==0 && local_vf_num==471 && local_vf_active==1) `fifo_error_check(471)
              else if (local_pf_num==0 && local_vf_num==472 && local_vf_active==1) `fifo_error_check(472)
              else if (local_pf_num==0 && local_vf_num==473 && local_vf_active==1) `fifo_error_check(473)
              else if (local_pf_num==0 && local_vf_num==474 && local_vf_active==1) `fifo_error_check(474)
              else if (local_pf_num==0 && local_vf_num==475 && local_vf_active==1) `fifo_error_check(475)
              else if (local_pf_num==0 && local_vf_num==476 && local_vf_active==1) `fifo_error_check(476)
              else if (local_pf_num==0 && local_vf_num==477 && local_vf_active==1) `fifo_error_check(477)
              else if (local_pf_num==0 && local_vf_num==478 && local_vf_active==1) `fifo_error_check(478)
              else if (local_pf_num==0 && local_vf_num==479 && local_vf_active==1) `fifo_error_check(479)
              else if (local_pf_num==0 && local_vf_num==480 && local_vf_active==1) `fifo_error_check(480)
              else if (local_pf_num==0 && local_vf_num==481 && local_vf_active==1) `fifo_error_check(481)
              else if (local_pf_num==0 && local_vf_num==482 && local_vf_active==1) `fifo_error_check(482)
              else if (local_pf_num==0 && local_vf_num==483 && local_vf_active==1) `fifo_error_check(483)
              else if (local_pf_num==0 && local_vf_num==484 && local_vf_active==1) `fifo_error_check(484)
              else if (local_pf_num==0 && local_vf_num==485 && local_vf_active==1) `fifo_error_check(485)
              else if (local_pf_num==0 && local_vf_num==486 && local_vf_active==1) `fifo_error_check(486)
              else if (local_pf_num==0 && local_vf_num==487 && local_vf_active==1) `fifo_error_check(487)
              else if (local_pf_num==0 && local_vf_num==488 && local_vf_active==1) `fifo_error_check(488)
              else if (local_pf_num==0 && local_vf_num==489 && local_vf_active==1) `fifo_error_check(489)
              else if (local_pf_num==0 && local_vf_num==490 && local_vf_active==1) `fifo_error_check(490)
              else if (local_pf_num==0 && local_vf_num==491 && local_vf_active==1) `fifo_error_check(491)
              else if (local_pf_num==0 && local_vf_num==492 && local_vf_active==1) `fifo_error_check(492)
              else if (local_pf_num==0 && local_vf_num==493 && local_vf_active==1) `fifo_error_check(493)
              else if (local_pf_num==0 && local_vf_num==494 && local_vf_active==1) `fifo_error_check(494)
              else if (local_pf_num==0 && local_vf_num==495 && local_vf_active==1) `fifo_error_check(495)
              else if (local_pf_num==0 && local_vf_num==496 && local_vf_active==1) `fifo_error_check(496)
              else if (local_pf_num==0 && local_vf_num==497 && local_vf_active==1) `fifo_error_check(497)
              else if (local_pf_num==0 && local_vf_num==498 && local_vf_active==1) `fifo_error_check(498)
              else if (local_pf_num==0 && local_vf_num==499 && local_vf_active==1) `fifo_error_check(499)
              else if (local_pf_num==0 && local_vf_num==500 && local_vf_active==1) `fifo_error_check(500)
              else if (local_pf_num==0 && local_vf_num==501 && local_vf_active==1) `fifo_error_check(501)
              else if (local_pf_num==0 && local_vf_num==502 && local_vf_active==1) `fifo_error_check(502)
              else if (local_pf_num==0 && local_vf_num==503 && local_vf_active==1) `fifo_error_check(503)
              else if (local_pf_num==0 && local_vf_num==504 && local_vf_active==1) `fifo_error_check(504)
              else if (local_pf_num==0 && local_vf_num==505 && local_vf_active==1) `fifo_error_check(505)
              else if (local_pf_num==0 && local_vf_num==506 && local_vf_active==1) `fifo_error_check(506)
              else if (local_pf_num==0 && local_vf_num==507 && local_vf_active==1) `fifo_error_check(507)
              else if (local_pf_num==0 && local_vf_num==508 && local_vf_active==1) `fifo_error_check(508)
              else if (local_pf_num==0 && local_vf_num==509 && local_vf_active==1) `fifo_error_check(509)
              else if (local_pf_num==0 && local_vf_num==510 && local_vf_active==1) `fifo_error_check(510)
              else if (local_pf_num==0 && local_vf_num==511 && local_vf_active==1) `fifo_error_check(511)
              else if (local_pf_num==0 && local_vf_num==512 && local_vf_active==1) `fifo_error_check(512)
              else if (local_pf_num==0 && local_vf_num==513 && local_vf_active==1) `fifo_error_check(513)
              else if (local_pf_num==0 && local_vf_num==514 && local_vf_active==1) `fifo_error_check(514)
              else if (local_pf_num==0 && local_vf_num==515 && local_vf_active==1) `fifo_error_check(515)
              else if (local_pf_num==0 && local_vf_num==516 && local_vf_active==1) `fifo_error_check(516)
              else if (local_pf_num==0 && local_vf_num==517 && local_vf_active==1) `fifo_error_check(517)
              else if (local_pf_num==0 && local_vf_num==518 && local_vf_active==1) `fifo_error_check(518)
              else if (local_pf_num==0 && local_vf_num==519 && local_vf_active==1) `fifo_error_check(519)
              else if (local_pf_num==0 && local_vf_num==520 && local_vf_active==1) `fifo_error_check(520)
              else if (local_pf_num==0 && local_vf_num==521 && local_vf_active==1) `fifo_error_check(521)
              else if (local_pf_num==0 && local_vf_num==522 && local_vf_active==1) `fifo_error_check(522)
              else if (local_pf_num==0 && local_vf_num==523 && local_vf_active==1) `fifo_error_check(523)
              else if (local_pf_num==0 && local_vf_num==524 && local_vf_active==1) `fifo_error_check(524)
              else if (local_pf_num==0 && local_vf_num==525 && local_vf_active==1) `fifo_error_check(525)
              else if (local_pf_num==0 && local_vf_num==526 && local_vf_active==1) `fifo_error_check(526)
              else if (local_pf_num==0 && local_vf_num==527 && local_vf_active==1) `fifo_error_check(527)
              else if (local_pf_num==0 && local_vf_num==528 && local_vf_active==1) `fifo_error_check(528)
              else if (local_pf_num==0 && local_vf_num==529 && local_vf_active==1) `fifo_error_check(529)
              else if (local_pf_num==0 && local_vf_num==530 && local_vf_active==1) `fifo_error_check(530)
              else if (local_pf_num==0 && local_vf_num==531 && local_vf_active==1) `fifo_error_check(531)
              else if (local_pf_num==0 && local_vf_num==532 && local_vf_active==1) `fifo_error_check(532)
              else if (local_pf_num==0 && local_vf_num==533 && local_vf_active==1) `fifo_error_check(533)
              else if (local_pf_num==0 && local_vf_num==534 && local_vf_active==1) `fifo_error_check(534)
              else if (local_pf_num==0 && local_vf_num==535 && local_vf_active==1) `fifo_error_check(535)
              else if (local_pf_num==0 && local_vf_num==536 && local_vf_active==1) `fifo_error_check(536)
              else if (local_pf_num==0 && local_vf_num==537 && local_vf_active==1) `fifo_error_check(537)
              else if (local_pf_num==0 && local_vf_num==538 && local_vf_active==1) `fifo_error_check(538)
              else if (local_pf_num==0 && local_vf_num==539 && local_vf_active==1) `fifo_error_check(539)
              else if (local_pf_num==0 && local_vf_num==540 && local_vf_active==1) `fifo_error_check(540)
              else if (local_pf_num==0 && local_vf_num==541 && local_vf_active==1) `fifo_error_check(541)
              else if (local_pf_num==0 && local_vf_num==542 && local_vf_active==1) `fifo_error_check(542)
              else if (local_pf_num==0 && local_vf_num==543 && local_vf_active==1) `fifo_error_check(543)
              else if (local_pf_num==0 && local_vf_num==544 && local_vf_active==1) `fifo_error_check(544)
              else if (local_pf_num==0 && local_vf_num==545 && local_vf_active==1) `fifo_error_check(545)
              else if (local_pf_num==0 && local_vf_num==546 && local_vf_active==1) `fifo_error_check(546)
              else if (local_pf_num==0 && local_vf_num==547 && local_vf_active==1) `fifo_error_check(547)
              else if (local_pf_num==0 && local_vf_num==548 && local_vf_active==1) `fifo_error_check(548)
              else if (local_pf_num==0 && local_vf_num==549 && local_vf_active==1) `fifo_error_check(549)
              else if (local_pf_num==0 && local_vf_num==550 && local_vf_active==1) `fifo_error_check(550)
              else if (local_pf_num==0 && local_vf_num==551 && local_vf_active==1) `fifo_error_check(551)
              else if (local_pf_num==0 && local_vf_num==552 && local_vf_active==1) `fifo_error_check(552)
              else if (local_pf_num==0 && local_vf_num==553 && local_vf_active==1) `fifo_error_check(553)
              else if (local_pf_num==0 && local_vf_num==554 && local_vf_active==1) `fifo_error_check(554)
              else if (local_pf_num==0 && local_vf_num==555 && local_vf_active==1) `fifo_error_check(555)
              else if (local_pf_num==0 && local_vf_num==556 && local_vf_active==1) `fifo_error_check(556)
              else if (local_pf_num==0 && local_vf_num==557 && local_vf_active==1) `fifo_error_check(557)
              else if (local_pf_num==0 && local_vf_num==558 && local_vf_active==1) `fifo_error_check(558)
              else if (local_pf_num==0 && local_vf_num==559 && local_vf_active==1) `fifo_error_check(559)
              else if (local_pf_num==0 && local_vf_num==560 && local_vf_active==1) `fifo_error_check(560)
              else if (local_pf_num==0 && local_vf_num==561 && local_vf_active==1) `fifo_error_check(561)
              else if (local_pf_num==0 && local_vf_num==562 && local_vf_active==1) `fifo_error_check(562)
              else if (local_pf_num==0 && local_vf_num==563 && local_vf_active==1) `fifo_error_check(563)
              else if (local_pf_num==0 && local_vf_num==564 && local_vf_active==1) `fifo_error_check(564)
              else if (local_pf_num==0 && local_vf_num==565 && local_vf_active==1) `fifo_error_check(565)
              else if (local_pf_num==0 && local_vf_num==566 && local_vf_active==1) `fifo_error_check(566)
              else if (local_pf_num==0 && local_vf_num==567 && local_vf_active==1) `fifo_error_check(567)
              else if (local_pf_num==0 && local_vf_num==568 && local_vf_active==1) `fifo_error_check(568)
              else if (local_pf_num==0 && local_vf_num==569 && local_vf_active==1) `fifo_error_check(569)
              else if (local_pf_num==0 && local_vf_num==570 && local_vf_active==1) `fifo_error_check(570)
              else if (local_pf_num==0 && local_vf_num==571 && local_vf_active==1) `fifo_error_check(571)
              else if (local_pf_num==0 && local_vf_num==572 && local_vf_active==1) `fifo_error_check(572)
              else if (local_pf_num==0 && local_vf_num==573 && local_vf_active==1) `fifo_error_check(573)
              else if (local_pf_num==0 && local_vf_num==574 && local_vf_active==1) `fifo_error_check(574)
              else if (local_pf_num==0 && local_vf_num==575 && local_vf_active==1) `fifo_error_check(575)
              else if (local_pf_num==0 && local_vf_num==576 && local_vf_active==1) `fifo_error_check(576)
              else if (local_pf_num==0 && local_vf_num==577 && local_vf_active==1) `fifo_error_check(577)
              else if (local_pf_num==0 && local_vf_num==578 && local_vf_active==1) `fifo_error_check(578)
              else if (local_pf_num==0 && local_vf_num==579 && local_vf_active==1) `fifo_error_check(579)
              else if (local_pf_num==0 && local_vf_num==580 && local_vf_active==1) `fifo_error_check(580)
              else if (local_pf_num==0 && local_vf_num==581 && local_vf_active==1) `fifo_error_check(581)
              else if (local_pf_num==0 && local_vf_num==582 && local_vf_active==1) `fifo_error_check(582)
              else if (local_pf_num==0 && local_vf_num==583 && local_vf_active==1) `fifo_error_check(583)
              else if (local_pf_num==0 && local_vf_num==584 && local_vf_active==1) `fifo_error_check(584)
              else if (local_pf_num==0 && local_vf_num==585 && local_vf_active==1) `fifo_error_check(585)
              else if (local_pf_num==0 && local_vf_num==586 && local_vf_active==1) `fifo_error_check(586)
              else if (local_pf_num==0 && local_vf_num==587 && local_vf_active==1) `fifo_error_check(587)
              else if (local_pf_num==0 && local_vf_num==588 && local_vf_active==1) `fifo_error_check(588)
              else if (local_pf_num==0 && local_vf_num==589 && local_vf_active==1) `fifo_error_check(589)
              else if (local_pf_num==0 && local_vf_num==590 && local_vf_active==1) `fifo_error_check(590)
              else if (local_pf_num==0 && local_vf_num==591 && local_vf_active==1) `fifo_error_check(591)
              else if (local_pf_num==0 && local_vf_num==592 && local_vf_active==1) `fifo_error_check(592)
              else if (local_pf_num==0 && local_vf_num==593 && local_vf_active==1) `fifo_error_check(593)
              else if (local_pf_num==0 && local_vf_num==594 && local_vf_active==1) `fifo_error_check(594)
              else if (local_pf_num==0 && local_vf_num==595 && local_vf_active==1) `fifo_error_check(595)
              else if (local_pf_num==0 && local_vf_num==596 && local_vf_active==1) `fifo_error_check(596)
              else if (local_pf_num==0 && local_vf_num==597 && local_vf_active==1) `fifo_error_check(597)
              else if (local_pf_num==0 && local_vf_num==598 && local_vf_active==1) `fifo_error_check(598)
              else if (local_pf_num==0 && local_vf_num==599 && local_vf_active==1) `fifo_error_check(599)
              else if (local_pf_num==0 && local_vf_num==600 && local_vf_active==1) `fifo_error_check(600)
              else if (local_pf_num==0 && local_vf_num==601 && local_vf_active==1) `fifo_error_check(601)
              else if (local_pf_num==0 && local_vf_num==602 && local_vf_active==1) `fifo_error_check(602)
              else if (local_pf_num==0 && local_vf_num==603 && local_vf_active==1) `fifo_error_check(603)
              else if (local_pf_num==0 && local_vf_num==604 && local_vf_active==1) `fifo_error_check(604)
              else if (local_pf_num==0 && local_vf_num==605 && local_vf_active==1) `fifo_error_check(605)
              else if (local_pf_num==0 && local_vf_num==606 && local_vf_active==1) `fifo_error_check(606)
              else if (local_pf_num==0 && local_vf_num==607 && local_vf_active==1) `fifo_error_check(607)
              else if (local_pf_num==0 && local_vf_num==608 && local_vf_active==1) `fifo_error_check(608)
              else if (local_pf_num==0 && local_vf_num==609 && local_vf_active==1) `fifo_error_check(609)
              else if (local_pf_num==0 && local_vf_num==610 && local_vf_active==1) `fifo_error_check(610)
              else if (local_pf_num==0 && local_vf_num==611 && local_vf_active==1) `fifo_error_check(611)
              else if (local_pf_num==0 && local_vf_num==612 && local_vf_active==1) `fifo_error_check(612)
              else if (local_pf_num==0 && local_vf_num==613 && local_vf_active==1) `fifo_error_check(613)
              else if (local_pf_num==0 && local_vf_num==614 && local_vf_active==1) `fifo_error_check(614)
              else if (local_pf_num==0 && local_vf_num==615 && local_vf_active==1) `fifo_error_check(615)
              else if (local_pf_num==0 && local_vf_num==616 && local_vf_active==1) `fifo_error_check(616)
              else if (local_pf_num==0 && local_vf_num==617 && local_vf_active==1) `fifo_error_check(617)
              else if (local_pf_num==0 && local_vf_num==618 && local_vf_active==1) `fifo_error_check(618)
              else if (local_pf_num==0 && local_vf_num==619 && local_vf_active==1) `fifo_error_check(619)
              else if (local_pf_num==0 && local_vf_num==620 && local_vf_active==1) `fifo_error_check(620)
              else if (local_pf_num==0 && local_vf_num==621 && local_vf_active==1) `fifo_error_check(621)
              else if (local_pf_num==0 && local_vf_num==622 && local_vf_active==1) `fifo_error_check(622)
              else if (local_pf_num==0 && local_vf_num==623 && local_vf_active==1) `fifo_error_check(623)
              else if (local_pf_num==0 && local_vf_num==624 && local_vf_active==1) `fifo_error_check(624)
              else if (local_pf_num==0 && local_vf_num==625 && local_vf_active==1) `fifo_error_check(625)
              else if (local_pf_num==0 && local_vf_num==626 && local_vf_active==1) `fifo_error_check(626)
              else if (local_pf_num==0 && local_vf_num==627 && local_vf_active==1) `fifo_error_check(627)
              else if (local_pf_num==0 && local_vf_num==628 && local_vf_active==1) `fifo_error_check(628)
              else if (local_pf_num==0 && local_vf_num==629 && local_vf_active==1) `fifo_error_check(629)
              else if (local_pf_num==0 && local_vf_num==630 && local_vf_active==1) `fifo_error_check(630)
              else if (local_pf_num==0 && local_vf_num==631 && local_vf_active==1) `fifo_error_check(631)
              else if (local_pf_num==0 && local_vf_num==632 && local_vf_active==1) `fifo_error_check(632)
              else if (local_pf_num==0 && local_vf_num==633 && local_vf_active==1) `fifo_error_check(633)
              else if (local_pf_num==0 && local_vf_num==634 && local_vf_active==1) `fifo_error_check(634)
              else if (local_pf_num==0 && local_vf_num==635 && local_vf_active==1) `fifo_error_check(635)
              else if (local_pf_num==0 && local_vf_num==636 && local_vf_active==1) `fifo_error_check(636)
              else if (local_pf_num==0 && local_vf_num==637 && local_vf_active==1) `fifo_error_check(637)
              else if (local_pf_num==0 && local_vf_num==638 && local_vf_active==1) `fifo_error_check(638)
              else if (local_pf_num==0 && local_vf_num==639 && local_vf_active==1) `fifo_error_check(639)
              else if (local_pf_num==0 && local_vf_num==640 && local_vf_active==1) `fifo_error_check(640)
              else if (local_pf_num==0 && local_vf_num==641 && local_vf_active==1) `fifo_error_check(641)
              else if (local_pf_num==0 && local_vf_num==642 && local_vf_active==1) `fifo_error_check(642)
              else if (local_pf_num==0 && local_vf_num==643 && local_vf_active==1) `fifo_error_check(643)
              else if (local_pf_num==0 && local_vf_num==644 && local_vf_active==1) `fifo_error_check(644)
              else if (local_pf_num==0 && local_vf_num==645 && local_vf_active==1) `fifo_error_check(645)
              else if (local_pf_num==0 && local_vf_num==646 && local_vf_active==1) `fifo_error_check(646)
              else if (local_pf_num==0 && local_vf_num==647 && local_vf_active==1) `fifo_error_check(647)
              else if (local_pf_num==0 && local_vf_num==648 && local_vf_active==1) `fifo_error_check(648)
              else if (local_pf_num==0 && local_vf_num==649 && local_vf_active==1) `fifo_error_check(649)
              else if (local_pf_num==0 && local_vf_num==650 && local_vf_active==1) `fifo_error_check(650)
              else if (local_pf_num==0 && local_vf_num==651 && local_vf_active==1) `fifo_error_check(651)
              else if (local_pf_num==0 && local_vf_num==652 && local_vf_active==1) `fifo_error_check(652)
              else if (local_pf_num==0 && local_vf_num==653 && local_vf_active==1) `fifo_error_check(653)
              else if (local_pf_num==0 && local_vf_num==654 && local_vf_active==1) `fifo_error_check(654)
              else if (local_pf_num==0 && local_vf_num==655 && local_vf_active==1) `fifo_error_check(655)
              else if (local_pf_num==0 && local_vf_num==656 && local_vf_active==1) `fifo_error_check(656)
              else if (local_pf_num==0 && local_vf_num==657 && local_vf_active==1) `fifo_error_check(657)
              else if (local_pf_num==0 && local_vf_num==658 && local_vf_active==1) `fifo_error_check(658)
              else if (local_pf_num==0 && local_vf_num==659 && local_vf_active==1) `fifo_error_check(659)
              else if (local_pf_num==0 && local_vf_num==660 && local_vf_active==1) `fifo_error_check(660)
              else if (local_pf_num==0 && local_vf_num==661 && local_vf_active==1) `fifo_error_check(661)
              else if (local_pf_num==0 && local_vf_num==662 && local_vf_active==1) `fifo_error_check(662)
              else if (local_pf_num==0 && local_vf_num==663 && local_vf_active==1) `fifo_error_check(663)
              else if (local_pf_num==0 && local_vf_num==664 && local_vf_active==1) `fifo_error_check(664)
              else if (local_pf_num==0 && local_vf_num==665 && local_vf_active==1) `fifo_error_check(665)
              else if (local_pf_num==0 && local_vf_num==666 && local_vf_active==1) `fifo_error_check(666)
              else if (local_pf_num==0 && local_vf_num==667 && local_vf_active==1) `fifo_error_check(667)
              else if (local_pf_num==0 && local_vf_num==668 && local_vf_active==1) `fifo_error_check(668)
              else if (local_pf_num==0 && local_vf_num==669 && local_vf_active==1) `fifo_error_check(669)
              else if (local_pf_num==0 && local_vf_num==670 && local_vf_active==1) `fifo_error_check(670)
              else if (local_pf_num==0 && local_vf_num==671 && local_vf_active==1) `fifo_error_check(671)
              else if (local_pf_num==0 && local_vf_num==672 && local_vf_active==1) `fifo_error_check(672)
              else if (local_pf_num==0 && local_vf_num==673 && local_vf_active==1) `fifo_error_check(673)
              else if (local_pf_num==0 && local_vf_num==674 && local_vf_active==1) `fifo_error_check(674)
              else if (local_pf_num==0 && local_vf_num==675 && local_vf_active==1) `fifo_error_check(675)
              else if (local_pf_num==0 && local_vf_num==676 && local_vf_active==1) `fifo_error_check(676)
              else if (local_pf_num==0 && local_vf_num==677 && local_vf_active==1) `fifo_error_check(677)
              else if (local_pf_num==0 && local_vf_num==678 && local_vf_active==1) `fifo_error_check(678)
              else if (local_pf_num==0 && local_vf_num==679 && local_vf_active==1) `fifo_error_check(679)
              else if (local_pf_num==0 && local_vf_num==680 && local_vf_active==1) `fifo_error_check(680)
              else if (local_pf_num==0 && local_vf_num==681 && local_vf_active==1) `fifo_error_check(681)
              else if (local_pf_num==0 && local_vf_num==682 && local_vf_active==1) `fifo_error_check(682)
              else if (local_pf_num==0 && local_vf_num==683 && local_vf_active==1) `fifo_error_check(683)
              else if (local_pf_num==0 && local_vf_num==684 && local_vf_active==1) `fifo_error_check(684)
              else if (local_pf_num==0 && local_vf_num==685 && local_vf_active==1) `fifo_error_check(685)
              else if (local_pf_num==0 && local_vf_num==686 && local_vf_active==1) `fifo_error_check(686)
              else if (local_pf_num==0 && local_vf_num==687 && local_vf_active==1) `fifo_error_check(687)
              else if (local_pf_num==0 && local_vf_num==688 && local_vf_active==1) `fifo_error_check(688)
              else if (local_pf_num==0 && local_vf_num==689 && local_vf_active==1) `fifo_error_check(689)
              else if (local_pf_num==0 && local_vf_num==690 && local_vf_active==1) `fifo_error_check(690)
              else if (local_pf_num==0 && local_vf_num==691 && local_vf_active==1) `fifo_error_check(691)
              else if (local_pf_num==0 && local_vf_num==692 && local_vf_active==1) `fifo_error_check(692)
              else if (local_pf_num==0 && local_vf_num==693 && local_vf_active==1) `fifo_error_check(693)
              else if (local_pf_num==0 && local_vf_num==694 && local_vf_active==1) `fifo_error_check(694)
              else if (local_pf_num==0 && local_vf_num==695 && local_vf_active==1) `fifo_error_check(695)
              else if (local_pf_num==0 && local_vf_num==696 && local_vf_active==1) `fifo_error_check(696)
              else if (local_pf_num==0 && local_vf_num==697 && local_vf_active==1) `fifo_error_check(697)
              else if (local_pf_num==0 && local_vf_num==698 && local_vf_active==1) `fifo_error_check(698)
              else if (local_pf_num==0 && local_vf_num==699 && local_vf_active==1) `fifo_error_check(699)
              else if (local_pf_num==0 && local_vf_num==700 && local_vf_active==1) `fifo_error_check(700)
              else if (local_pf_num==0 && local_vf_num==701 && local_vf_active==1) `fifo_error_check(701)
              else if (local_pf_num==0 && local_vf_num==702 && local_vf_active==1) `fifo_error_check(702)
              else if (local_pf_num==0 && local_vf_num==703 && local_vf_active==1) `fifo_error_check(703)
              else if (local_pf_num==0 && local_vf_num==704 && local_vf_active==1) `fifo_error_check(704)
              else if (local_pf_num==0 && local_vf_num==705 && local_vf_active==1) `fifo_error_check(705)
              else if (local_pf_num==0 && local_vf_num==706 && local_vf_active==1) `fifo_error_check(706)
              else if (local_pf_num==0 && local_vf_num==707 && local_vf_active==1) `fifo_error_check(707)
              else if (local_pf_num==0 && local_vf_num==708 && local_vf_active==1) `fifo_error_check(708)
              else if (local_pf_num==0 && local_vf_num==709 && local_vf_active==1) `fifo_error_check(709)
              else if (local_pf_num==0 && local_vf_num==710 && local_vf_active==1) `fifo_error_check(710)
              else if (local_pf_num==0 && local_vf_num==711 && local_vf_active==1) `fifo_error_check(711)
              else if (local_pf_num==0 && local_vf_num==712 && local_vf_active==1) `fifo_error_check(712)
              else if (local_pf_num==0 && local_vf_num==713 && local_vf_active==1) `fifo_error_check(713)
              else if (local_pf_num==0 && local_vf_num==714 && local_vf_active==1) `fifo_error_check(714)
              else if (local_pf_num==0 && local_vf_num==715 && local_vf_active==1) `fifo_error_check(715)
              else if (local_pf_num==0 && local_vf_num==716 && local_vf_active==1) `fifo_error_check(716)
              else if (local_pf_num==0 && local_vf_num==717 && local_vf_active==1) `fifo_error_check(717)
              else if (local_pf_num==0 && local_vf_num==718 && local_vf_active==1) `fifo_error_check(718)
              else if (local_pf_num==0 && local_vf_num==719 && local_vf_active==1) `fifo_error_check(719)
              else if (local_pf_num==0 && local_vf_num==720 && local_vf_active==1) `fifo_error_check(720)
              else if (local_pf_num==0 && local_vf_num==721 && local_vf_active==1) `fifo_error_check(721)
              else if (local_pf_num==0 && local_vf_num==722 && local_vf_active==1) `fifo_error_check(722)
              else if (local_pf_num==0 && local_vf_num==723 && local_vf_active==1) `fifo_error_check(723)
              else if (local_pf_num==0 && local_vf_num==724 && local_vf_active==1) `fifo_error_check(724)
              else if (local_pf_num==0 && local_vf_num==725 && local_vf_active==1) `fifo_error_check(725)
              else if (local_pf_num==0 && local_vf_num==726 && local_vf_active==1) `fifo_error_check(726)
              else if (local_pf_num==0 && local_vf_num==727 && local_vf_active==1) `fifo_error_check(727)
              else if (local_pf_num==0 && local_vf_num==728 && local_vf_active==1) `fifo_error_check(728)
              else if (local_pf_num==0 && local_vf_num==729 && local_vf_active==1) `fifo_error_check(729)
              else if (local_pf_num==0 && local_vf_num==730 && local_vf_active==1) `fifo_error_check(730)
              else if (local_pf_num==0 && local_vf_num==731 && local_vf_active==1) `fifo_error_check(731)
              else if (local_pf_num==0 && local_vf_num==732 && local_vf_active==1) `fifo_error_check(732)
              else if (local_pf_num==0 && local_vf_num==733 && local_vf_active==1) `fifo_error_check(733)
              else if (local_pf_num==0 && local_vf_num==734 && local_vf_active==1) `fifo_error_check(734)
              else if (local_pf_num==0 && local_vf_num==735 && local_vf_active==1) `fifo_error_check(735)
              else if (local_pf_num==0 && local_vf_num==736 && local_vf_active==1) `fifo_error_check(736)
              else if (local_pf_num==0 && local_vf_num==737 && local_vf_active==1) `fifo_error_check(737)
              else if (local_pf_num==0 && local_vf_num==738 && local_vf_active==1) `fifo_error_check(738)
              else if (local_pf_num==0 && local_vf_num==739 && local_vf_active==1) `fifo_error_check(739)
              else if (local_pf_num==0 && local_vf_num==740 && local_vf_active==1) `fifo_error_check(740)
              else if (local_pf_num==0 && local_vf_num==741 && local_vf_active==1) `fifo_error_check(741)
              else if (local_pf_num==0 && local_vf_num==742 && local_vf_active==1) `fifo_error_check(742)
              else if (local_pf_num==0 && local_vf_num==743 && local_vf_active==1) `fifo_error_check(743)
              else if (local_pf_num==0 && local_vf_num==744 && local_vf_active==1) `fifo_error_check(744)
              else if (local_pf_num==0 && local_vf_num==745 && local_vf_active==1) `fifo_error_check(745)
              else if (local_pf_num==0 && local_vf_num==746 && local_vf_active==1) `fifo_error_check(746)
              else if (local_pf_num==0 && local_vf_num==747 && local_vf_active==1) `fifo_error_check(747)
              else if (local_pf_num==0 && local_vf_num==748 && local_vf_active==1) `fifo_error_check(748)
              else if (local_pf_num==0 && local_vf_num==749 && local_vf_active==1) `fifo_error_check(749)
              else if (local_pf_num==0 && local_vf_num==750 && local_vf_active==1) `fifo_error_check(750)
              else if (local_pf_num==0 && local_vf_num==751 && local_vf_active==1) `fifo_error_check(751)
              else if (local_pf_num==0 && local_vf_num==752 && local_vf_active==1) `fifo_error_check(752)
              else if (local_pf_num==0 && local_vf_num==753 && local_vf_active==1) `fifo_error_check(753)
              else if (local_pf_num==0 && local_vf_num==754 && local_vf_active==1) `fifo_error_check(754)
              else if (local_pf_num==0 && local_vf_num==755 && local_vf_active==1) `fifo_error_check(755)
              else if (local_pf_num==0 && local_vf_num==756 && local_vf_active==1) `fifo_error_check(756)
              else if (local_pf_num==0 && local_vf_num==757 && local_vf_active==1) `fifo_error_check(757)
              else if (local_pf_num==0 && local_vf_num==758 && local_vf_active==1) `fifo_error_check(758)
              else if (local_pf_num==0 && local_vf_num==759 && local_vf_active==1) `fifo_error_check(759)
              else if (local_pf_num==0 && local_vf_num==760 && local_vf_active==1) `fifo_error_check(760)
              else if (local_pf_num==0 && local_vf_num==761 && local_vf_active==1) `fifo_error_check(761)
              else if (local_pf_num==0 && local_vf_num==762 && local_vf_active==1) `fifo_error_check(762)
              else if (local_pf_num==0 && local_vf_num==763 && local_vf_active==1) `fifo_error_check(763)
              else if (local_pf_num==0 && local_vf_num==764 && local_vf_active==1) `fifo_error_check(764)
              else if (local_pf_num==0 && local_vf_num==765 && local_vf_active==1) `fifo_error_check(765)
              else if (local_pf_num==0 && local_vf_num==766 && local_vf_active==1) `fifo_error_check(766)
              else if (local_pf_num==0 && local_vf_num==767 && local_vf_active==1) `fifo_error_check(767)
              else if (local_pf_num==0 && local_vf_num==768 && local_vf_active==1) `fifo_error_check(768)
              else if (local_pf_num==0 && local_vf_num==769 && local_vf_active==1) `fifo_error_check(769)
              else if (local_pf_num==0 && local_vf_num==770 && local_vf_active==1) `fifo_error_check(770)
              else if (local_pf_num==0 && local_vf_num==771 && local_vf_active==1) `fifo_error_check(771)
              else if (local_pf_num==0 && local_vf_num==772 && local_vf_active==1) `fifo_error_check(772)
              else if (local_pf_num==0 && local_vf_num==773 && local_vf_active==1) `fifo_error_check(773)
              else if (local_pf_num==0 && local_vf_num==774 && local_vf_active==1) `fifo_error_check(774)
              else if (local_pf_num==0 && local_vf_num==775 && local_vf_active==1) `fifo_error_check(775)
              else if (local_pf_num==0 && local_vf_num==776 && local_vf_active==1) `fifo_error_check(776)
              else if (local_pf_num==0 && local_vf_num==777 && local_vf_active==1) `fifo_error_check(777)
              else if (local_pf_num==0 && local_vf_num==778 && local_vf_active==1) `fifo_error_check(778)
              else if (local_pf_num==0 && local_vf_num==779 && local_vf_active==1) `fifo_error_check(779)
              else if (local_pf_num==0 && local_vf_num==780 && local_vf_active==1) `fifo_error_check(780)
              else if (local_pf_num==0 && local_vf_num==781 && local_vf_active==1) `fifo_error_check(781)
              else if (local_pf_num==0 && local_vf_num==782 && local_vf_active==1) `fifo_error_check(782)
              else if (local_pf_num==0 && local_vf_num==783 && local_vf_active==1) `fifo_error_check(783)
              else if (local_pf_num==0 && local_vf_num==784 && local_vf_active==1) `fifo_error_check(784)
              else if (local_pf_num==0 && local_vf_num==785 && local_vf_active==1) `fifo_error_check(785)
              else if (local_pf_num==0 && local_vf_num==786 && local_vf_active==1) `fifo_error_check(786)
              else if (local_pf_num==0 && local_vf_num==787 && local_vf_active==1) `fifo_error_check(787)
              else if (local_pf_num==0 && local_vf_num==788 && local_vf_active==1) `fifo_error_check(788)
              else if (local_pf_num==0 && local_vf_num==789 && local_vf_active==1) `fifo_error_check(789)
              else if (local_pf_num==0 && local_vf_num==790 && local_vf_active==1) `fifo_error_check(790)
              else if (local_pf_num==0 && local_vf_num==791 && local_vf_active==1) `fifo_error_check(791)
              else if (local_pf_num==0 && local_vf_num==792 && local_vf_active==1) `fifo_error_check(792)
              else if (local_pf_num==0 && local_vf_num==793 && local_vf_active==1) `fifo_error_check(793)
              else if (local_pf_num==0 && local_vf_num==794 && local_vf_active==1) `fifo_error_check(794)
              else if (local_pf_num==0 && local_vf_num==795 && local_vf_active==1) `fifo_error_check(795)
              else if (local_pf_num==0 && local_vf_num==796 && local_vf_active==1) `fifo_error_check(796)
              else if (local_pf_num==0 && local_vf_num==797 && local_vf_active==1) `fifo_error_check(797)
              else if (local_pf_num==0 && local_vf_num==798 && local_vf_active==1) `fifo_error_check(798)
              else if (local_pf_num==0 && local_vf_num==799 && local_vf_active==1) `fifo_error_check(799)
              else if (local_pf_num==0 && local_vf_num==800 && local_vf_active==1) `fifo_error_check(800)
              else if (local_pf_num==0 && local_vf_num==801 && local_vf_active==1) `fifo_error_check(801)
              else if (local_pf_num==0 && local_vf_num==802 && local_vf_active==1) `fifo_error_check(802)
              else if (local_pf_num==0 && local_vf_num==803 && local_vf_active==1) `fifo_error_check(803)
              else if (local_pf_num==0 && local_vf_num==804 && local_vf_active==1) `fifo_error_check(804)
              else if (local_pf_num==0 && local_vf_num==805 && local_vf_active==1) `fifo_error_check(805)
              else if (local_pf_num==0 && local_vf_num==806 && local_vf_active==1) `fifo_error_check(806)
              else if (local_pf_num==0 && local_vf_num==807 && local_vf_active==1) `fifo_error_check(807)
              else if (local_pf_num==0 && local_vf_num==808 && local_vf_active==1) `fifo_error_check(808)
              else if (local_pf_num==0 && local_vf_num==809 && local_vf_active==1) `fifo_error_check(809)
              else if (local_pf_num==0 && local_vf_num==810 && local_vf_active==1) `fifo_error_check(810)
              else if (local_pf_num==0 && local_vf_num==811 && local_vf_active==1) `fifo_error_check(811)
              else if (local_pf_num==0 && local_vf_num==812 && local_vf_active==1) `fifo_error_check(812)
              else if (local_pf_num==0 && local_vf_num==813 && local_vf_active==1) `fifo_error_check(813)
              else if (local_pf_num==0 && local_vf_num==814 && local_vf_active==1) `fifo_error_check(814)
              else if (local_pf_num==0 && local_vf_num==815 && local_vf_active==1) `fifo_error_check(815)
              else if (local_pf_num==0 && local_vf_num==816 && local_vf_active==1) `fifo_error_check(816)
              else if (local_pf_num==0 && local_vf_num==817 && local_vf_active==1) `fifo_error_check(817)
              else if (local_pf_num==0 && local_vf_num==818 && local_vf_active==1) `fifo_error_check(818)
              else if (local_pf_num==0 && local_vf_num==819 && local_vf_active==1) `fifo_error_check(819)
              else if (local_pf_num==0 && local_vf_num==820 && local_vf_active==1) `fifo_error_check(820)
              else if (local_pf_num==0 && local_vf_num==821 && local_vf_active==1) `fifo_error_check(821)
              else if (local_pf_num==0 && local_vf_num==822 && local_vf_active==1) `fifo_error_check(822)
              else if (local_pf_num==0 && local_vf_num==823 && local_vf_active==1) `fifo_error_check(823)
              else if (local_pf_num==0 && local_vf_num==824 && local_vf_active==1) `fifo_error_check(824)
              else if (local_pf_num==0 && local_vf_num==825 && local_vf_active==1) `fifo_error_check(825)
              else if (local_pf_num==0 && local_vf_num==826 && local_vf_active==1) `fifo_error_check(826)
              else if (local_pf_num==0 && local_vf_num==827 && local_vf_active==1) `fifo_error_check(827)
              else if (local_pf_num==0 && local_vf_num==828 && local_vf_active==1) `fifo_error_check(828)
              else if (local_pf_num==0 && local_vf_num==829 && local_vf_active==1) `fifo_error_check(829)
              else if (local_pf_num==0 && local_vf_num==830 && local_vf_active==1) `fifo_error_check(830)
              else if (local_pf_num==0 && local_vf_num==831 && local_vf_active==1) `fifo_error_check(831)
              else if (local_pf_num==0 && local_vf_num==832 && local_vf_active==1) `fifo_error_check(832)
              else if (local_pf_num==0 && local_vf_num==833 && local_vf_active==1) `fifo_error_check(833)
              else if (local_pf_num==0 && local_vf_num==834 && local_vf_active==1) `fifo_error_check(834)
              else if (local_pf_num==0 && local_vf_num==835 && local_vf_active==1) `fifo_error_check(835)
              else if (local_pf_num==0 && local_vf_num==836 && local_vf_active==1) `fifo_error_check(836)
              else if (local_pf_num==0 && local_vf_num==837 && local_vf_active==1) `fifo_error_check(837)
              else if (local_pf_num==0 && local_vf_num==838 && local_vf_active==1) `fifo_error_check(838)
              else if (local_pf_num==0 && local_vf_num==839 && local_vf_active==1) `fifo_error_check(839)
              else if (local_pf_num==0 && local_vf_num==840 && local_vf_active==1) `fifo_error_check(840)
              else if (local_pf_num==0 && local_vf_num==841 && local_vf_active==1) `fifo_error_check(841)
              else if (local_pf_num==0 && local_vf_num==842 && local_vf_active==1) `fifo_error_check(842)
              else if (local_pf_num==0 && local_vf_num==843 && local_vf_active==1) `fifo_error_check(843)
              else if (local_pf_num==0 && local_vf_num==844 && local_vf_active==1) `fifo_error_check(844)
              else if (local_pf_num==0 && local_vf_num==845 && local_vf_active==1) `fifo_error_check(845)
              else if (local_pf_num==0 && local_vf_num==846 && local_vf_active==1) `fifo_error_check(846)
              else if (local_pf_num==0 && local_vf_num==847 && local_vf_active==1) `fifo_error_check(847)
              else if (local_pf_num==0 && local_vf_num==848 && local_vf_active==1) `fifo_error_check(848)
              else if (local_pf_num==0 && local_vf_num==849 && local_vf_active==1) `fifo_error_check(849)
              else if (local_pf_num==0 && local_vf_num==850 && local_vf_active==1) `fifo_error_check(850)
              else if (local_pf_num==0 && local_vf_num==851 && local_vf_active==1) `fifo_error_check(851)
              else if (local_pf_num==0 && local_vf_num==852 && local_vf_active==1) `fifo_error_check(852)
              else if (local_pf_num==0 && local_vf_num==853 && local_vf_active==1) `fifo_error_check(853)
              else if (local_pf_num==0 && local_vf_num==854 && local_vf_active==1) `fifo_error_check(854)
              else if (local_pf_num==0 && local_vf_num==855 && local_vf_active==1) `fifo_error_check(855)
              else if (local_pf_num==0 && local_vf_num==856 && local_vf_active==1) `fifo_error_check(856)
              else if (local_pf_num==0 && local_vf_num==857 && local_vf_active==1) `fifo_error_check(857)
              else if (local_pf_num==0 && local_vf_num==858 && local_vf_active==1) `fifo_error_check(858)
              else if (local_pf_num==0 && local_vf_num==859 && local_vf_active==1) `fifo_error_check(859)
              else if (local_pf_num==0 && local_vf_num==860 && local_vf_active==1) `fifo_error_check(860)
              else if (local_pf_num==0 && local_vf_num==861 && local_vf_active==1) `fifo_error_check(861)
              else if (local_pf_num==0 && local_vf_num==862 && local_vf_active==1) `fifo_error_check(862)
              else if (local_pf_num==0 && local_vf_num==863 && local_vf_active==1) `fifo_error_check(863)
              else if (local_pf_num==0 && local_vf_num==864 && local_vf_active==1) `fifo_error_check(864)
              else if (local_pf_num==0 && local_vf_num==865 && local_vf_active==1) `fifo_error_check(865)
              else if (local_pf_num==0 && local_vf_num==866 && local_vf_active==1) `fifo_error_check(866)
              else if (local_pf_num==0 && local_vf_num==867 && local_vf_active==1) `fifo_error_check(867)
              else if (local_pf_num==0 && local_vf_num==868 && local_vf_active==1) `fifo_error_check(868)
              else if (local_pf_num==0 && local_vf_num==869 && local_vf_active==1) `fifo_error_check(869)
              else if (local_pf_num==0 && local_vf_num==870 && local_vf_active==1) `fifo_error_check(870)
              else if (local_pf_num==0 && local_vf_num==871 && local_vf_active==1) `fifo_error_check(871)
              else if (local_pf_num==0 && local_vf_num==872 && local_vf_active==1) `fifo_error_check(872)
              else if (local_pf_num==0 && local_vf_num==873 && local_vf_active==1) `fifo_error_check(873)
              else if (local_pf_num==0 && local_vf_num==874 && local_vf_active==1) `fifo_error_check(874)
              else if (local_pf_num==0 && local_vf_num==875 && local_vf_active==1) `fifo_error_check(875)
              else if (local_pf_num==0 && local_vf_num==876 && local_vf_active==1) `fifo_error_check(876)
              else if (local_pf_num==0 && local_vf_num==877 && local_vf_active==1) `fifo_error_check(877)
              else if (local_pf_num==0 && local_vf_num==878 && local_vf_active==1) `fifo_error_check(878)
              else if (local_pf_num==0 && local_vf_num==879 && local_vf_active==1) `fifo_error_check(879)
              else if (local_pf_num==0 && local_vf_num==880 && local_vf_active==1) `fifo_error_check(880)
              else if (local_pf_num==0 && local_vf_num==881 && local_vf_active==1) `fifo_error_check(881)
              else if (local_pf_num==0 && local_vf_num==882 && local_vf_active==1) `fifo_error_check(882)
              else if (local_pf_num==0 && local_vf_num==883 && local_vf_active==1) `fifo_error_check(883)
              else if (local_pf_num==0 && local_vf_num==884 && local_vf_active==1) `fifo_error_check(884)
              else if (local_pf_num==0 && local_vf_num==885 && local_vf_active==1) `fifo_error_check(885)
              else if (local_pf_num==0 && local_vf_num==886 && local_vf_active==1) `fifo_error_check(886)
              else if (local_pf_num==0 && local_vf_num==887 && local_vf_active==1) `fifo_error_check(887)
              else if (local_pf_num==0 && local_vf_num==888 && local_vf_active==1) `fifo_error_check(888)
              else if (local_pf_num==0 && local_vf_num==889 && local_vf_active==1) `fifo_error_check(889)
              else if (local_pf_num==0 && local_vf_num==890 && local_vf_active==1) `fifo_error_check(890)
              else if (local_pf_num==0 && local_vf_num==891 && local_vf_active==1) `fifo_error_check(891)
              else if (local_pf_num==0 && local_vf_num==892 && local_vf_active==1) `fifo_error_check(892)
              else if (local_pf_num==0 && local_vf_num==893 && local_vf_active==1) `fifo_error_check(893)
              else if (local_pf_num==0 && local_vf_num==894 && local_vf_active==1) `fifo_error_check(894)
              else if (local_pf_num==0 && local_vf_num==895 && local_vf_active==1) `fifo_error_check(895)
              else if (local_pf_num==0 && local_vf_num==896 && local_vf_active==1) `fifo_error_check(896)
              else if (local_pf_num==0 && local_vf_num==897 && local_vf_active==1) `fifo_error_check(897)
              else if (local_pf_num==0 && local_vf_num==898 && local_vf_active==1) `fifo_error_check(898)
              else if (local_pf_num==0 && local_vf_num==899 && local_vf_active==1) `fifo_error_check(899)
              else if (local_pf_num==0 && local_vf_num==900 && local_vf_active==1) `fifo_error_check(900)
              else if (local_pf_num==0 && local_vf_num==901 && local_vf_active==1) `fifo_error_check(901)
              else if (local_pf_num==0 && local_vf_num==902 && local_vf_active==1) `fifo_error_check(902)
              else if (local_pf_num==0 && local_vf_num==903 && local_vf_active==1) `fifo_error_check(903)
              else if (local_pf_num==0 && local_vf_num==904 && local_vf_active==1) `fifo_error_check(904)
              else if (local_pf_num==0 && local_vf_num==905 && local_vf_active==1) `fifo_error_check(905)
              else if (local_pf_num==0 && local_vf_num==906 && local_vf_active==1) `fifo_error_check(906)
              else if (local_pf_num==0 && local_vf_num==907 && local_vf_active==1) `fifo_error_check(907)
              else if (local_pf_num==0 && local_vf_num==908 && local_vf_active==1) `fifo_error_check(908)
              else if (local_pf_num==0 && local_vf_num==909 && local_vf_active==1) `fifo_error_check(909)
              else if (local_pf_num==0 && local_vf_num==910 && local_vf_active==1) `fifo_error_check(910)
              else if (local_pf_num==0 && local_vf_num==911 && local_vf_active==1) `fifo_error_check(911)
              else if (local_pf_num==0 && local_vf_num==912 && local_vf_active==1) `fifo_error_check(912)
              else if (local_pf_num==0 && local_vf_num==913 && local_vf_active==1) `fifo_error_check(913)
              else if (local_pf_num==0 && local_vf_num==914 && local_vf_active==1) `fifo_error_check(914)
              else if (local_pf_num==0 && local_vf_num==915 && local_vf_active==1) `fifo_error_check(915)
              else if (local_pf_num==0 && local_vf_num==916 && local_vf_active==1) `fifo_error_check(916)
              else if (local_pf_num==0 && local_vf_num==917 && local_vf_active==1) `fifo_error_check(917)
              else if (local_pf_num==0 && local_vf_num==918 && local_vf_active==1) `fifo_error_check(918)
              else if (local_pf_num==0 && local_vf_num==919 && local_vf_active==1) `fifo_error_check(919)
              else if (local_pf_num==0 && local_vf_num==920 && local_vf_active==1) `fifo_error_check(920)
              else if (local_pf_num==0 && local_vf_num==921 && local_vf_active==1) `fifo_error_check(921)
              else if (local_pf_num==0 && local_vf_num==922 && local_vf_active==1) `fifo_error_check(922)
              else if (local_pf_num==0 && local_vf_num==923 && local_vf_active==1) `fifo_error_check(923)
              else if (local_pf_num==0 && local_vf_num==924 && local_vf_active==1) `fifo_error_check(924)
              else if (local_pf_num==0 && local_vf_num==925 && local_vf_active==1) `fifo_error_check(925)
              else if (local_pf_num==0 && local_vf_num==926 && local_vf_active==1) `fifo_error_check(926)
              else if (local_pf_num==0 && local_vf_num==927 && local_vf_active==1) `fifo_error_check(927)
              else if (local_pf_num==0 && local_vf_num==928 && local_vf_active==1) `fifo_error_check(928)
              else if (local_pf_num==0 && local_vf_num==929 && local_vf_active==1) `fifo_error_check(929)
              else if (local_pf_num==0 && local_vf_num==930 && local_vf_active==1) `fifo_error_check(930)
              else if (local_pf_num==0 && local_vf_num==931 && local_vf_active==1) `fifo_error_check(931)
              else if (local_pf_num==0 && local_vf_num==932 && local_vf_active==1) `fifo_error_check(932)
              else if (local_pf_num==0 && local_vf_num==933 && local_vf_active==1) `fifo_error_check(933)
              else if (local_pf_num==0 && local_vf_num==934 && local_vf_active==1) `fifo_error_check(934)
              else if (local_pf_num==0 && local_vf_num==935 && local_vf_active==1) `fifo_error_check(935)
              else if (local_pf_num==0 && local_vf_num==936 && local_vf_active==1) `fifo_error_check(936)
              else if (local_pf_num==0 && local_vf_num==937 && local_vf_active==1) `fifo_error_check(937)
              else if (local_pf_num==0 && local_vf_num==938 && local_vf_active==1) `fifo_error_check(938)
              else if (local_pf_num==0 && local_vf_num==939 && local_vf_active==1) `fifo_error_check(939)
              else if (local_pf_num==0 && local_vf_num==940 && local_vf_active==1) `fifo_error_check(940)
              else if (local_pf_num==0 && local_vf_num==941 && local_vf_active==1) `fifo_error_check(941)
              else if (local_pf_num==0 && local_vf_num==942 && local_vf_active==1) `fifo_error_check(942)
              else if (local_pf_num==0 && local_vf_num==943 && local_vf_active==1) `fifo_error_check(943)
              else if (local_pf_num==0 && local_vf_num==944 && local_vf_active==1) `fifo_error_check(944)
              else if (local_pf_num==0 && local_vf_num==945 && local_vf_active==1) `fifo_error_check(945)
              else if (local_pf_num==0 && local_vf_num==946 && local_vf_active==1) `fifo_error_check(946)
              else if (local_pf_num==0 && local_vf_num==947 && local_vf_active==1) `fifo_error_check(947)
              else if (local_pf_num==0 && local_vf_num==948 && local_vf_active==1) `fifo_error_check(948)
              else if (local_pf_num==0 && local_vf_num==949 && local_vf_active==1) `fifo_error_check(949)
              else if (local_pf_num==0 && local_vf_num==950 && local_vf_active==1) `fifo_error_check(950)
              else if (local_pf_num==0 && local_vf_num==951 && local_vf_active==1) `fifo_error_check(951)
              else if (local_pf_num==0 && local_vf_num==952 && local_vf_active==1) `fifo_error_check(952)
              else if (local_pf_num==0 && local_vf_num==953 && local_vf_active==1) `fifo_error_check(953)
              else if (local_pf_num==0 && local_vf_num==954 && local_vf_active==1) `fifo_error_check(954)
              else if (local_pf_num==0 && local_vf_num==955 && local_vf_active==1) `fifo_error_check(955)
              else if (local_pf_num==0 && local_vf_num==956 && local_vf_active==1) `fifo_error_check(956)
              else if (local_pf_num==0 && local_vf_num==957 && local_vf_active==1) `fifo_error_check(957)
              else if (local_pf_num==0 && local_vf_num==958 && local_vf_active==1) `fifo_error_check(958)
              else if (local_pf_num==0 && local_vf_num==959 && local_vf_active==1) `fifo_error_check(959)
              else if (local_pf_num==0 && local_vf_num==960 && local_vf_active==1) `fifo_error_check(960)
              else if (local_pf_num==0 && local_vf_num==961 && local_vf_active==1) `fifo_error_check(961)
              else if (local_pf_num==0 && local_vf_num==962 && local_vf_active==1) `fifo_error_check(962)
              else if (local_pf_num==0 && local_vf_num==963 && local_vf_active==1) `fifo_error_check(963)
              else if (local_pf_num==0 && local_vf_num==964 && local_vf_active==1) `fifo_error_check(964)
              else if (local_pf_num==0 && local_vf_num==965 && local_vf_active==1) `fifo_error_check(965)
              else if (local_pf_num==0 && local_vf_num==966 && local_vf_active==1) `fifo_error_check(966)
              else if (local_pf_num==0 && local_vf_num==967 && local_vf_active==1) `fifo_error_check(967)
              else if (local_pf_num==0 && local_vf_num==968 && local_vf_active==1) `fifo_error_check(968)
              else if (local_pf_num==0 && local_vf_num==969 && local_vf_active==1) `fifo_error_check(969)
              else if (local_pf_num==0 && local_vf_num==970 && local_vf_active==1) `fifo_error_check(970)
              else if (local_pf_num==0 && local_vf_num==971 && local_vf_active==1) `fifo_error_check(971)
              else if (local_pf_num==0 && local_vf_num==972 && local_vf_active==1) `fifo_error_check(972)
              else if (local_pf_num==0 && local_vf_num==973 && local_vf_active==1) `fifo_error_check(973)
              else if (local_pf_num==0 && local_vf_num==974 && local_vf_active==1) `fifo_error_check(974)
              else if (local_pf_num==0 && local_vf_num==975 && local_vf_active==1) `fifo_error_check(975)
              else if (local_pf_num==0 && local_vf_num==976 && local_vf_active==1) `fifo_error_check(976)
              else if (local_pf_num==0 && local_vf_num==977 && local_vf_active==1) `fifo_error_check(977)
              else if (local_pf_num==0 && local_vf_num==978 && local_vf_active==1) `fifo_error_check(978)
              else if (local_pf_num==0 && local_vf_num==979 && local_vf_active==1) `fifo_error_check(979)
              else if (local_pf_num==0 && local_vf_num==980 && local_vf_active==1) `fifo_error_check(980)
              else if (local_pf_num==0 && local_vf_num==981 && local_vf_active==1) `fifo_error_check(981)
              else if (local_pf_num==0 && local_vf_num==982 && local_vf_active==1) `fifo_error_check(982)
              else if (local_pf_num==0 && local_vf_num==983 && local_vf_active==1) `fifo_error_check(983)
              else if (local_pf_num==0 && local_vf_num==984 && local_vf_active==1) `fifo_error_check(984)
              else if (local_pf_num==0 && local_vf_num==985 && local_vf_active==1) `fifo_error_check(985)
              else if (local_pf_num==0 && local_vf_num==986 && local_vf_active==1) `fifo_error_check(986)
              else if (local_pf_num==0 && local_vf_num==987 && local_vf_active==1) `fifo_error_check(987)
              else if (local_pf_num==0 && local_vf_num==988 && local_vf_active==1) `fifo_error_check(988)
              else if (local_pf_num==0 && local_vf_num==989 && local_vf_active==1) `fifo_error_check(989)
              else if (local_pf_num==0 && local_vf_num==990 && local_vf_active==1) `fifo_error_check(990)
              else if (local_pf_num==0 && local_vf_num==991 && local_vf_active==1) `fifo_error_check(991)
              else if (local_pf_num==0 && local_vf_num==992 && local_vf_active==1) `fifo_error_check(992)
              else if (local_pf_num==0 && local_vf_num==993 && local_vf_active==1) `fifo_error_check(993)
              else if (local_pf_num==0 && local_vf_num==994 && local_vf_active==1) `fifo_error_check(994)
              else if (local_pf_num==0 && local_vf_num==995 && local_vf_active==1) `fifo_error_check(995)
              else if (local_pf_num==0 && local_vf_num==996 && local_vf_active==1) `fifo_error_check(996)
              else if (local_pf_num==0 && local_vf_num==997 && local_vf_active==1) `fifo_error_check(997)
              else if (local_pf_num==0 && local_vf_num==998 && local_vf_active==1) `fifo_error_check(998)
              else if (local_pf_num==0 && local_vf_num==999 && local_vf_active==1) `fifo_error_check(999)
              else if (local_pf_num==0 && local_vf_num==1000 && local_vf_active==1) `fifo_error_check(1000)
              else if (local_pf_num==0 && local_vf_num==1001 && local_vf_active==1) `fifo_error_check(1001)
              else if (local_pf_num==0 && local_vf_num==1002 && local_vf_active==1) `fifo_error_check(1002)
              else if (local_pf_num==0 && local_vf_num==1003 && local_vf_active==1) `fifo_error_check(1003)
              else if (local_pf_num==0 && local_vf_num==1004 && local_vf_active==1) `fifo_error_check(1004)
              else if (local_pf_num==0 && local_vf_num==1005 && local_vf_active==1) `fifo_error_check(1005)
              else if (local_pf_num==0 && local_vf_num==1006 && local_vf_active==1) `fifo_error_check(1006)
              else if (local_pf_num==0 && local_vf_num==1007 && local_vf_active==1) `fifo_error_check(1007)
              else if (local_pf_num==0 && local_vf_num==1008 && local_vf_active==1) `fifo_error_check(1008)
              else if (local_pf_num==0 && local_vf_num==1009 && local_vf_active==1) `fifo_error_check(1009)
              else if (local_pf_num==0 && local_vf_num==1010 && local_vf_active==1) `fifo_error_check(1010)
              else if (local_pf_num==0 && local_vf_num==1011 && local_vf_active==1) `fifo_error_check(1011)
              else if (local_pf_num==0 && local_vf_num==1012 && local_vf_active==1) `fifo_error_check(1012)
              else if (local_pf_num==0 && local_vf_num==1013 && local_vf_active==1) `fifo_error_check(1013)
              else if (local_pf_num==0 && local_vf_num==1014 && local_vf_active==1) `fifo_error_check(1014)
              else if (local_pf_num==0 && local_vf_num==1015 && local_vf_active==1) `fifo_error_check(1015)
              else if (local_pf_num==0 && local_vf_num==1016 && local_vf_active==1) `fifo_error_check(1016)
              else if (local_pf_num==0 && local_vf_num==1017 && local_vf_active==1) `fifo_error_check(1017)
              else if (local_pf_num==0 && local_vf_num==1018 && local_vf_active==1) `fifo_error_check(1018)
              else if (local_pf_num==0 && local_vf_num==1019 && local_vf_active==1) `fifo_error_check(1019)
              else if (local_pf_num==0 && local_vf_num==1020 && local_vf_active==1) `fifo_error_check(1020)
              else if (local_pf_num==0 && local_vf_num==1021 && local_vf_active==1) `fifo_error_check(1021)
              else if (local_pf_num==0 && local_vf_num==1022 && local_vf_active==1) `fifo_error_check(1022)
              else if (local_pf_num==0 && local_vf_num==1023 && local_vf_active==1) `fifo_error_check(1023)
              else if (local_pf_num==0 && local_vf_num==1024 && local_vf_active==1) `fifo_error_check(1024)
              else if (local_pf_num==0 && local_vf_num==1025 && local_vf_active==1) `fifo_error_check(1025)
              else if (local_pf_num==0 && local_vf_num==1026 && local_vf_active==1) `fifo_error_check(1026)
              else if (local_pf_num==0 && local_vf_num==1027 && local_vf_active==1) `fifo_error_check(1027)
              else if (local_pf_num==0 && local_vf_num==1028 && local_vf_active==1) `fifo_error_check(1028)
              else if (local_pf_num==0 && local_vf_num==1029 && local_vf_active==1) `fifo_error_check(1029)
              else if (local_pf_num==0 && local_vf_num==1030 && local_vf_active==1) `fifo_error_check(1030)
              else if (local_pf_num==0 && local_vf_num==1031 && local_vf_active==1) `fifo_error_check(1031)
              else if (local_pf_num==0 && local_vf_num==1032 && local_vf_active==1) `fifo_error_check(1032)
              else if (local_pf_num==0 && local_vf_num==1033 && local_vf_active==1) `fifo_error_check(1033)
              else if (local_pf_num==0 && local_vf_num==1034 && local_vf_active==1) `fifo_error_check(1034)
              else if (local_pf_num==0 && local_vf_num==1035 && local_vf_active==1) `fifo_error_check(1035)
              else if (local_pf_num==0 && local_vf_num==1036 && local_vf_active==1) `fifo_error_check(1036)
              else if (local_pf_num==0 && local_vf_num==1037 && local_vf_active==1) `fifo_error_check(1037)
              else if (local_pf_num==0 && local_vf_num==1038 && local_vf_active==1) `fifo_error_check(1038)
              else if (local_pf_num==0 && local_vf_num==1039 && local_vf_active==1) `fifo_error_check(1039)
              else if (local_pf_num==0 && local_vf_num==1040 && local_vf_active==1) `fifo_error_check(1040)
              else if (local_pf_num==0 && local_vf_num==1041 && local_vf_active==1) `fifo_error_check(1041)
              else if (local_pf_num==0 && local_vf_num==1042 && local_vf_active==1) `fifo_error_check(1042)
              else if (local_pf_num==0 && local_vf_num==1043 && local_vf_active==1) `fifo_error_check(1043)
              else if (local_pf_num==0 && local_vf_num==1044 && local_vf_active==1) `fifo_error_check(1044)
              else if (local_pf_num==0 && local_vf_num==1045 && local_vf_active==1) `fifo_error_check(1045)
              else if (local_pf_num==0 && local_vf_num==1046 && local_vf_active==1) `fifo_error_check(1046)
              else if (local_pf_num==0 && local_vf_num==1047 && local_vf_active==1) `fifo_error_check(1047)
              else if (local_pf_num==0 && local_vf_num==1048 && local_vf_active==1) `fifo_error_check(1048)
              else if (local_pf_num==0 && local_vf_num==1049 && local_vf_active==1) `fifo_error_check(1049)
              else if (local_pf_num==0 && local_vf_num==1050 && local_vf_active==1) `fifo_error_check(1050)
              else if (local_pf_num==0 && local_vf_num==1051 && local_vf_active==1) `fifo_error_check(1051)
              else if (local_pf_num==0 && local_vf_num==1052 && local_vf_active==1) `fifo_error_check(1052)
              else if (local_pf_num==0 && local_vf_num==1053 && local_vf_active==1) `fifo_error_check(1053)
              else if (local_pf_num==0 && local_vf_num==1054 && local_vf_active==1) `fifo_error_check(1054)
              else if (local_pf_num==0 && local_vf_num==1055 && local_vf_active==1) `fifo_error_check(1055)
              else if (local_pf_num==0 && local_vf_num==1056 && local_vf_active==1) `fifo_error_check(1056)
              else if (local_pf_num==0 && local_vf_num==1057 && local_vf_active==1) `fifo_error_check(1057)
              else if (local_pf_num==0 && local_vf_num==1058 && local_vf_active==1) `fifo_error_check(1058)
              else if (local_pf_num==0 && local_vf_num==1059 && local_vf_active==1) `fifo_error_check(1059)
              else if (local_pf_num==0 && local_vf_num==1060 && local_vf_active==1) `fifo_error_check(1060)
              else if (local_pf_num==0 && local_vf_num==1061 && local_vf_active==1) `fifo_error_check(1061)
              else if (local_pf_num==0 && local_vf_num==1062 && local_vf_active==1) `fifo_error_check(1062)
              else if (local_pf_num==0 && local_vf_num==1063 && local_vf_active==1) `fifo_error_check(1063)
              else if (local_pf_num==0 && local_vf_num==1064 && local_vf_active==1) `fifo_error_check(1064)
              else if (local_pf_num==0 && local_vf_num==1065 && local_vf_active==1) `fifo_error_check(1065)
              else if (local_pf_num==0 && local_vf_num==1066 && local_vf_active==1) `fifo_error_check(1066)
              else if (local_pf_num==0 && local_vf_num==1067 && local_vf_active==1) `fifo_error_check(1067)
              else if (local_pf_num==0 && local_vf_num==1068 && local_vf_active==1) `fifo_error_check(1068)
              else if (local_pf_num==0 && local_vf_num==1069 && local_vf_active==1) `fifo_error_check(1069)
              else if (local_pf_num==0 && local_vf_num==1070 && local_vf_active==1) `fifo_error_check(1070)
              else if (local_pf_num==0 && local_vf_num==1071 && local_vf_active==1) `fifo_error_check(1071)
              else if (local_pf_num==0 && local_vf_num==1072 && local_vf_active==1) `fifo_error_check(1072)
              else if (local_pf_num==0 && local_vf_num==1073 && local_vf_active==1) `fifo_error_check(1073)
              else if (local_pf_num==0 && local_vf_num==1074 && local_vf_active==1) `fifo_error_check(1074)
              else if (local_pf_num==0 && local_vf_num==1075 && local_vf_active==1) `fifo_error_check(1075)
              else if (local_pf_num==0 && local_vf_num==1076 && local_vf_active==1) `fifo_error_check(1076)
              else if (local_pf_num==0 && local_vf_num==1077 && local_vf_active==1) `fifo_error_check(1077)
              else if (local_pf_num==0 && local_vf_num==1078 && local_vf_active==1) `fifo_error_check(1078)
              else if (local_pf_num==0 && local_vf_num==1079 && local_vf_active==1) `fifo_error_check(1079)
              else if (local_pf_num==0 && local_vf_num==1080 && local_vf_active==1) `fifo_error_check(1080)
              else if (local_pf_num==0 && local_vf_num==1081 && local_vf_active==1) `fifo_error_check(1081)
              else if (local_pf_num==0 && local_vf_num==1082 && local_vf_active==1) `fifo_error_check(1082)
              else if (local_pf_num==0 && local_vf_num==1083 && local_vf_active==1) `fifo_error_check(1083)
              else if (local_pf_num==0 && local_vf_num==1084 && local_vf_active==1) `fifo_error_check(1084)
              else if (local_pf_num==0 && local_vf_num==1085 && local_vf_active==1) `fifo_error_check(1085)
              else if (local_pf_num==0 && local_vf_num==1086 && local_vf_active==1) `fifo_error_check(1086)
              else if (local_pf_num==0 && local_vf_num==1087 && local_vf_active==1) `fifo_error_check(1087)
              else if (local_pf_num==0 && local_vf_num==1088 && local_vf_active==1) `fifo_error_check(1088)
              else if (local_pf_num==0 && local_vf_num==1089 && local_vf_active==1) `fifo_error_check(1089)
              else if (local_pf_num==0 && local_vf_num==1090 && local_vf_active==1) `fifo_error_check(1090)
              else if (local_pf_num==0 && local_vf_num==1091 && local_vf_active==1) `fifo_error_check(1091)
              else if (local_pf_num==0 && local_vf_num==1092 && local_vf_active==1) `fifo_error_check(1092)
              else if (local_pf_num==0 && local_vf_num==1093 && local_vf_active==1) `fifo_error_check(1093)
              else if (local_pf_num==0 && local_vf_num==1094 && local_vf_active==1) `fifo_error_check(1094)
              else if (local_pf_num==0 && local_vf_num==1095 && local_vf_active==1) `fifo_error_check(1095)
              else if (local_pf_num==0 && local_vf_num==1096 && local_vf_active==1) `fifo_error_check(1096)
              else if (local_pf_num==0 && local_vf_num==1097 && local_vf_active==1) `fifo_error_check(1097)
              else if (local_pf_num==0 && local_vf_num==1098 && local_vf_active==1) `fifo_error_check(1098)
              else if (local_pf_num==0 && local_vf_num==1099 && local_vf_active==1) `fifo_error_check(1099)
              else if (local_pf_num==0 && local_vf_num==1100 && local_vf_active==1) `fifo_error_check(1100)
              else if (local_pf_num==0 && local_vf_num==1101 && local_vf_active==1) `fifo_error_check(1101)
              else if (local_pf_num==0 && local_vf_num==1102 && local_vf_active==1) `fifo_error_check(1102)
              else if (local_pf_num==0 && local_vf_num==1103 && local_vf_active==1) `fifo_error_check(1103)
              else if (local_pf_num==0 && local_vf_num==1104 && local_vf_active==1) `fifo_error_check(1104)
              else if (local_pf_num==0 && local_vf_num==1105 && local_vf_active==1) `fifo_error_check(1105)
              else if (local_pf_num==0 && local_vf_num==1106 && local_vf_active==1) `fifo_error_check(1106)
              else if (local_pf_num==0 && local_vf_num==1107 && local_vf_active==1) `fifo_error_check(1107)
              else if (local_pf_num==0 && local_vf_num==1108 && local_vf_active==1) `fifo_error_check(1108)
              else if (local_pf_num==0 && local_vf_num==1109 && local_vf_active==1) `fifo_error_check(1109)
              else if (local_pf_num==0 && local_vf_num==1110 && local_vf_active==1) `fifo_error_check(1110)
              else if (local_pf_num==0 && local_vf_num==1111 && local_vf_active==1) `fifo_error_check(1111)
              else if (local_pf_num==0 && local_vf_num==1112 && local_vf_active==1) `fifo_error_check(1112)
              else if (local_pf_num==0 && local_vf_num==1113 && local_vf_active==1) `fifo_error_check(1113)
              else if (local_pf_num==0 && local_vf_num==1114 && local_vf_active==1) `fifo_error_check(1114)
              else if (local_pf_num==0 && local_vf_num==1115 && local_vf_active==1) `fifo_error_check(1115)
              else if (local_pf_num==0 && local_vf_num==1116 && local_vf_active==1) `fifo_error_check(1116)
              else if (local_pf_num==0 && local_vf_num==1117 && local_vf_active==1) `fifo_error_check(1117)
              else if (local_pf_num==0 && local_vf_num==1118 && local_vf_active==1) `fifo_error_check(1118)
              else if (local_pf_num==0 && local_vf_num==1119 && local_vf_active==1) `fifo_error_check(1119)
              else if (local_pf_num==0 && local_vf_num==1120 && local_vf_active==1) `fifo_error_check(1120)
              else if (local_pf_num==0 && local_vf_num==1121 && local_vf_active==1) `fifo_error_check(1121)
              else if (local_pf_num==0 && local_vf_num==1122 && local_vf_active==1) `fifo_error_check(1122)
              else if (local_pf_num==0 && local_vf_num==1123 && local_vf_active==1) `fifo_error_check(1123)
              else if (local_pf_num==0 && local_vf_num==1124 && local_vf_active==1) `fifo_error_check(1124)
              else if (local_pf_num==0 && local_vf_num==1125 && local_vf_active==1) `fifo_error_check(1125)
              else if (local_pf_num==0 && local_vf_num==1126 && local_vf_active==1) `fifo_error_check(1126)
              else if (local_pf_num==0 && local_vf_num==1127 && local_vf_active==1) `fifo_error_check(1127)
              else if (local_pf_num==0 && local_vf_num==1128 && local_vf_active==1) `fifo_error_check(1128)
              else if (local_pf_num==0 && local_vf_num==1129 && local_vf_active==1) `fifo_error_check(1129)
              else if (local_pf_num==0 && local_vf_num==1130 && local_vf_active==1) `fifo_error_check(1130)
              else if (local_pf_num==0 && local_vf_num==1131 && local_vf_active==1) `fifo_error_check(1131)
              else if (local_pf_num==0 && local_vf_num==1132 && local_vf_active==1) `fifo_error_check(1132)
              else if (local_pf_num==0 && local_vf_num==1133 && local_vf_active==1) `fifo_error_check(1133)
              else if (local_pf_num==0 && local_vf_num==1134 && local_vf_active==1) `fifo_error_check(1134)
              else if (local_pf_num==0 && local_vf_num==1135 && local_vf_active==1) `fifo_error_check(1135)
              else if (local_pf_num==0 && local_vf_num==1136 && local_vf_active==1) `fifo_error_check(1136)
              else if (local_pf_num==0 && local_vf_num==1137 && local_vf_active==1) `fifo_error_check(1137)
              else if (local_pf_num==0 && local_vf_num==1138 && local_vf_active==1) `fifo_error_check(1138)
              else if (local_pf_num==0 && local_vf_num==1139 && local_vf_active==1) `fifo_error_check(1139)
              else if (local_pf_num==0 && local_vf_num==1140 && local_vf_active==1) `fifo_error_check(1140)
              else if (local_pf_num==0 && local_vf_num==1141 && local_vf_active==1) `fifo_error_check(1141)
              else if (local_pf_num==0 && local_vf_num==1142 && local_vf_active==1) `fifo_error_check(1142)
              else if (local_pf_num==0 && local_vf_num==1143 && local_vf_active==1) `fifo_error_check(1143)
              else if (local_pf_num==0 && local_vf_num==1144 && local_vf_active==1) `fifo_error_check(1144)
              else if (local_pf_num==0 && local_vf_num==1145 && local_vf_active==1) `fifo_error_check(1145)
              else if (local_pf_num==0 && local_vf_num==1146 && local_vf_active==1) `fifo_error_check(1146)
              else if (local_pf_num==0 && local_vf_num==1147 && local_vf_active==1) `fifo_error_check(1147)
              else if (local_pf_num==0 && local_vf_num==1148 && local_vf_active==1) `fifo_error_check(1148)
              else if (local_pf_num==0 && local_vf_num==1149 && local_vf_active==1) `fifo_error_check(1149)
              else if (local_pf_num==0 && local_vf_num==1150 && local_vf_active==1) `fifo_error_check(1150)
              else if (local_pf_num==0 && local_vf_num==1151 && local_vf_active==1) `fifo_error_check(1151)
              else if (local_pf_num==0 && local_vf_num==1152 && local_vf_active==1) `fifo_error_check(1152)
              else if (local_pf_num==0 && local_vf_num==1153 && local_vf_active==1) `fifo_error_check(1153)
              else if (local_pf_num==0 && local_vf_num==1154 && local_vf_active==1) `fifo_error_check(1154)
              else if (local_pf_num==0 && local_vf_num==1155 && local_vf_active==1) `fifo_error_check(1155)
              else if (local_pf_num==0 && local_vf_num==1156 && local_vf_active==1) `fifo_error_check(1156)
              else if (local_pf_num==0 && local_vf_num==1157 && local_vf_active==1) `fifo_error_check(1157)
              else if (local_pf_num==0 && local_vf_num==1158 && local_vf_active==1) `fifo_error_check(1158)
              else if (local_pf_num==0 && local_vf_num==1159 && local_vf_active==1) `fifo_error_check(1159)
              else if (local_pf_num==0 && local_vf_num==1160 && local_vf_active==1) `fifo_error_check(1160)
              else if (local_pf_num==0 && local_vf_num==1161 && local_vf_active==1) `fifo_error_check(1161)
              else if (local_pf_num==0 && local_vf_num==1162 && local_vf_active==1) `fifo_error_check(1162)
              else if (local_pf_num==0 && local_vf_num==1163 && local_vf_active==1) `fifo_error_check(1163)
              else if (local_pf_num==0 && local_vf_num==1164 && local_vf_active==1) `fifo_error_check(1164)
              else if (local_pf_num==0 && local_vf_num==1165 && local_vf_active==1) `fifo_error_check(1165)
              else if (local_pf_num==0 && local_vf_num==1166 && local_vf_active==1) `fifo_error_check(1166)
              else if (local_pf_num==0 && local_vf_num==1167 && local_vf_active==1) `fifo_error_check(1167)
              else if (local_pf_num==0 && local_vf_num==1168 && local_vf_active==1) `fifo_error_check(1168)
              else if (local_pf_num==0 && local_vf_num==1169 && local_vf_active==1) `fifo_error_check(1169)
              else if (local_pf_num==0 && local_vf_num==1170 && local_vf_active==1) `fifo_error_check(1170)
              else if (local_pf_num==0 && local_vf_num==1171 && local_vf_active==1) `fifo_error_check(1171)
              else if (local_pf_num==0 && local_vf_num==1172 && local_vf_active==1) `fifo_error_check(1172)
              else if (local_pf_num==0 && local_vf_num==1173 && local_vf_active==1) `fifo_error_check(1173)
              else if (local_pf_num==0 && local_vf_num==1174 && local_vf_active==1) `fifo_error_check(1174)
              else if (local_pf_num==0 && local_vf_num==1175 && local_vf_active==1) `fifo_error_check(1175)
              else if (local_pf_num==0 && local_vf_num==1176 && local_vf_active==1) `fifo_error_check(1176)
              else if (local_pf_num==0 && local_vf_num==1177 && local_vf_active==1) `fifo_error_check(1177)
              else if (local_pf_num==0 && local_vf_num==1178 && local_vf_active==1) `fifo_error_check(1178)
              else if (local_pf_num==0 && local_vf_num==1179 && local_vf_active==1) `fifo_error_check(1179)
              else if (local_pf_num==0 && local_vf_num==1180 && local_vf_active==1) `fifo_error_check(1180)
              else if (local_pf_num==0 && local_vf_num==1181 && local_vf_active==1) `fifo_error_check(1181)
              else if (local_pf_num==0 && local_vf_num==1182 && local_vf_active==1) `fifo_error_check(1182)
              else if (local_pf_num==0 && local_vf_num==1183 && local_vf_active==1) `fifo_error_check(1183)
              else if (local_pf_num==0 && local_vf_num==1184 && local_vf_active==1) `fifo_error_check(1184)
              else if (local_pf_num==0 && local_vf_num==1185 && local_vf_active==1) `fifo_error_check(1185)
              else if (local_pf_num==0 && local_vf_num==1186 && local_vf_active==1) `fifo_error_check(1186)
              else if (local_pf_num==0 && local_vf_num==1187 && local_vf_active==1) `fifo_error_check(1187)
              else if (local_pf_num==0 && local_vf_num==1188 && local_vf_active==1) `fifo_error_check(1188)
              else if (local_pf_num==0 && local_vf_num==1189 && local_vf_active==1) `fifo_error_check(1189)
              else if (local_pf_num==0 && local_vf_num==1190 && local_vf_active==1) `fifo_error_check(1190)
              else if (local_pf_num==0 && local_vf_num==1191 && local_vf_active==1) `fifo_error_check(1191)
              else if (local_pf_num==0 && local_vf_num==1192 && local_vf_active==1) `fifo_error_check(1192)
              else if (local_pf_num==0 && local_vf_num==1193 && local_vf_active==1) `fifo_error_check(1193)
              else if (local_pf_num==0 && local_vf_num==1194 && local_vf_active==1) `fifo_error_check(1194)
              else if (local_pf_num==0 && local_vf_num==1195 && local_vf_active==1) `fifo_error_check(1195)
              else if (local_pf_num==0 && local_vf_num==1196 && local_vf_active==1) `fifo_error_check(1196)
              else if (local_pf_num==0 && local_vf_num==1197 && local_vf_active==1) `fifo_error_check(1197)
              else if (local_pf_num==0 && local_vf_num==1198 && local_vf_active==1) `fifo_error_check(1198)
              else if (local_pf_num==0 && local_vf_num==1199 && local_vf_active==1) `fifo_error_check(1199)
              else if (local_pf_num==0 && local_vf_num==1200 && local_vf_active==1) `fifo_error_check(1200)
              else if (local_pf_num==0 && local_vf_num==1201 && local_vf_active==1) `fifo_error_check(1201)
              else if (local_pf_num==0 && local_vf_num==1202 && local_vf_active==1) `fifo_error_check(1202)
              else if (local_pf_num==0 && local_vf_num==1203 && local_vf_active==1) `fifo_error_check(1203)
              else if (local_pf_num==0 && local_vf_num==1204 && local_vf_active==1) `fifo_error_check(1204)
              else if (local_pf_num==0 && local_vf_num==1205 && local_vf_active==1) `fifo_error_check(1205)
              else if (local_pf_num==0 && local_vf_num==1206 && local_vf_active==1) `fifo_error_check(1206)
              else if (local_pf_num==0 && local_vf_num==1207 && local_vf_active==1) `fifo_error_check(1207)
              else if (local_pf_num==0 && local_vf_num==1208 && local_vf_active==1) `fifo_error_check(1208)
              else if (local_pf_num==0 && local_vf_num==1209 && local_vf_active==1) `fifo_error_check(1209)
              else if (local_pf_num==0 && local_vf_num==1210 && local_vf_active==1) `fifo_error_check(1210)
              else if (local_pf_num==0 && local_vf_num==1211 && local_vf_active==1) `fifo_error_check(1211)
              else if (local_pf_num==0 && local_vf_num==1212 && local_vf_active==1) `fifo_error_check(1212)
              else if (local_pf_num==0 && local_vf_num==1213 && local_vf_active==1) `fifo_error_check(1213)
              else if (local_pf_num==0 && local_vf_num==1214 && local_vf_active==1) `fifo_error_check(1214)
              else if (local_pf_num==0 && local_vf_num==1215 && local_vf_active==1) `fifo_error_check(1215)
              else if (local_pf_num==0 && local_vf_num==1216 && local_vf_active==1) `fifo_error_check(1216)
              else if (local_pf_num==0 && local_vf_num==1217 && local_vf_active==1) `fifo_error_check(1217)
              else if (local_pf_num==0 && local_vf_num==1218 && local_vf_active==1) `fifo_error_check(1218)
              else if (local_pf_num==0 && local_vf_num==1219 && local_vf_active==1) `fifo_error_check(1219)
              else if (local_pf_num==0 && local_vf_num==1220 && local_vf_active==1) `fifo_error_check(1220)
              else if (local_pf_num==0 && local_vf_num==1221 && local_vf_active==1) `fifo_error_check(1221)
              else if (local_pf_num==0 && local_vf_num==1222 && local_vf_active==1) `fifo_error_check(1222)
              else if (local_pf_num==0 && local_vf_num==1223 && local_vf_active==1) `fifo_error_check(1223)
              else if (local_pf_num==0 && local_vf_num==1224 && local_vf_active==1) `fifo_error_check(1224)
              else if (local_pf_num==0 && local_vf_num==1225 && local_vf_active==1) `fifo_error_check(1225)
              else if (local_pf_num==0 && local_vf_num==1226 && local_vf_active==1) `fifo_error_check(1226)
              else if (local_pf_num==0 && local_vf_num==1227 && local_vf_active==1) `fifo_error_check(1227)
              else if (local_pf_num==0 && local_vf_num==1228 && local_vf_active==1) `fifo_error_check(1228)
              else if (local_pf_num==0 && local_vf_num==1229 && local_vf_active==1) `fifo_error_check(1229)
              else if (local_pf_num==0 && local_vf_num==1230 && local_vf_active==1) `fifo_error_check(1230)
              else if (local_pf_num==0 && local_vf_num==1231 && local_vf_active==1) `fifo_error_check(1231)
              else if (local_pf_num==0 && local_vf_num==1232 && local_vf_active==1) `fifo_error_check(1232)
              else if (local_pf_num==0 && local_vf_num==1233 && local_vf_active==1) `fifo_error_check(1233)
              else if (local_pf_num==0 && local_vf_num==1234 && local_vf_active==1) `fifo_error_check(1234)
              else if (local_pf_num==0 && local_vf_num==1235 && local_vf_active==1) `fifo_error_check(1235)
              else if (local_pf_num==0 && local_vf_num==1236 && local_vf_active==1) `fifo_error_check(1236)
              else if (local_pf_num==0 && local_vf_num==1237 && local_vf_active==1) `fifo_error_check(1237)
              else if (local_pf_num==0 && local_vf_num==1238 && local_vf_active==1) `fifo_error_check(1238)
              else if (local_pf_num==0 && local_vf_num==1239 && local_vf_active==1) `fifo_error_check(1239)
              else if (local_pf_num==0 && local_vf_num==1240 && local_vf_active==1) `fifo_error_check(1240)
              else if (local_pf_num==0 && local_vf_num==1241 && local_vf_active==1) `fifo_error_check(1241)
              else if (local_pf_num==0 && local_vf_num==1242 && local_vf_active==1) `fifo_error_check(1242)
              else if (local_pf_num==0 && local_vf_num==1243 && local_vf_active==1) `fifo_error_check(1243)
              else if (local_pf_num==0 && local_vf_num==1244 && local_vf_active==1) `fifo_error_check(1244)
              else if (local_pf_num==0 && local_vf_num==1245 && local_vf_active==1) `fifo_error_check(1245)
              else if (local_pf_num==0 && local_vf_num==1246 && local_vf_active==1) `fifo_error_check(1246)
              else if (local_pf_num==0 && local_vf_num==1247 && local_vf_active==1) `fifo_error_check(1247)
              else if (local_pf_num==0 && local_vf_num==1248 && local_vf_active==1) `fifo_error_check(1248)
              else if (local_pf_num==0 && local_vf_num==1249 && local_vf_active==1) `fifo_error_check(1249)
              else if (local_pf_num==0 && local_vf_num==1250 && local_vf_active==1) `fifo_error_check(1250)
              else if (local_pf_num==0 && local_vf_num==1251 && local_vf_active==1) `fifo_error_check(1251)
              else if (local_pf_num==0 && local_vf_num==1252 && local_vf_active==1) `fifo_error_check(1252)
              else if (local_pf_num==0 && local_vf_num==1253 && local_vf_active==1) `fifo_error_check(1253)
              else if (local_pf_num==0 && local_vf_num==1254 && local_vf_active==1) `fifo_error_check(1254)
              else if (local_pf_num==0 && local_vf_num==1255 && local_vf_active==1) `fifo_error_check(1255)
              else if (local_pf_num==0 && local_vf_num==1256 && local_vf_active==1) `fifo_error_check(1256)
              else if (local_pf_num==0 && local_vf_num==1257 && local_vf_active==1) `fifo_error_check(1257)
              else if (local_pf_num==0 && local_vf_num==1258 && local_vf_active==1) `fifo_error_check(1258)
              else if (local_pf_num==0 && local_vf_num==1259 && local_vf_active==1) `fifo_error_check(1259)
              else if (local_pf_num==0 && local_vf_num==1260 && local_vf_active==1) `fifo_error_check(1260)
              else if (local_pf_num==0 && local_vf_num==1261 && local_vf_active==1) `fifo_error_check(1261)
              else if (local_pf_num==0 && local_vf_num==1262 && local_vf_active==1) `fifo_error_check(1262)
              else if (local_pf_num==0 && local_vf_num==1263 && local_vf_active==1) `fifo_error_check(1263)
              else if (local_pf_num==0 && local_vf_num==1264 && local_vf_active==1) `fifo_error_check(1264)
              else if (local_pf_num==0 && local_vf_num==1265 && local_vf_active==1) `fifo_error_check(1265)
              else if (local_pf_num==0 && local_vf_num==1266 && local_vf_active==1) `fifo_error_check(1266)
              else if (local_pf_num==0 && local_vf_num==1267 && local_vf_active==1) `fifo_error_check(1267)
              else if (local_pf_num==0 && local_vf_num==1268 && local_vf_active==1) `fifo_error_check(1268)
              else if (local_pf_num==0 && local_vf_num==1269 && local_vf_active==1) `fifo_error_check(1269)
              else if (local_pf_num==0 && local_vf_num==1270 && local_vf_active==1) `fifo_error_check(1270)
              else if (local_pf_num==0 && local_vf_num==1271 && local_vf_active==1) `fifo_error_check(1271)
              else if (local_pf_num==0 && local_vf_num==1272 && local_vf_active==1) `fifo_error_check(1272)
              else if (local_pf_num==0 && local_vf_num==1273 && local_vf_active==1) `fifo_error_check(1273)
              else if (local_pf_num==0 && local_vf_num==1274 && local_vf_active==1) `fifo_error_check(1274)
              else if (local_pf_num==0 && local_vf_num==1275 && local_vf_active==1) `fifo_error_check(1275)
              else if (local_pf_num==0 && local_vf_num==1276 && local_vf_active==1) `fifo_error_check(1276)
              else if (local_pf_num==0 && local_vf_num==1277 && local_vf_active==1) `fifo_error_check(1277)
              else if (local_pf_num==0 && local_vf_num==1278 && local_vf_active==1) `fifo_error_check(1278)
              else if (local_pf_num==0 && local_vf_num==1279 && local_vf_active==1) `fifo_error_check(1279)
              else if (local_pf_num==0 && local_vf_num==1280 && local_vf_active==1) `fifo_error_check(1280)
              else if (local_pf_num==0 && local_vf_num==1281 && local_vf_active==1) `fifo_error_check(1281)
              else if (local_pf_num==0 && local_vf_num==1282 && local_vf_active==1) `fifo_error_check(1282)
              else if (local_pf_num==0 && local_vf_num==1283 && local_vf_active==1) `fifo_error_check(1283)
              else if (local_pf_num==0 && local_vf_num==1284 && local_vf_active==1) `fifo_error_check(1284)
              else if (local_pf_num==0 && local_vf_num==1285 && local_vf_active==1) `fifo_error_check(1285)
              else if (local_pf_num==0 && local_vf_num==1286 && local_vf_active==1) `fifo_error_check(1286)
              else if (local_pf_num==0 && local_vf_num==1287 && local_vf_active==1) `fifo_error_check(1287)
              else if (local_pf_num==0 && local_vf_num==1288 && local_vf_active==1) `fifo_error_check(1288)
              else if (local_pf_num==0 && local_vf_num==1289 && local_vf_active==1) `fifo_error_check(1289)
              else if (local_pf_num==0 && local_vf_num==1290 && local_vf_active==1) `fifo_error_check(1290)
              else if (local_pf_num==0 && local_vf_num==1291 && local_vf_active==1) `fifo_error_check(1291)
              else if (local_pf_num==0 && local_vf_num==1292 && local_vf_active==1) `fifo_error_check(1292)
              else if (local_pf_num==0 && local_vf_num==1293 && local_vf_active==1) `fifo_error_check(1293)
              else if (local_pf_num==0 && local_vf_num==1294 && local_vf_active==1) `fifo_error_check(1294)
              else if (local_pf_num==0 && local_vf_num==1295 && local_vf_active==1) `fifo_error_check(1295)
              else if (local_pf_num==0 && local_vf_num==1296 && local_vf_active==1) `fifo_error_check(1296)
              else if (local_pf_num==0 && local_vf_num==1297 && local_vf_active==1) `fifo_error_check(1297)
              else if (local_pf_num==0 && local_vf_num==1298 && local_vf_active==1) `fifo_error_check(1298)
              else if (local_pf_num==0 && local_vf_num==1299 && local_vf_active==1) `fifo_error_check(1299)
              else if (local_pf_num==0 && local_vf_num==1300 && local_vf_active==1) `fifo_error_check(1300)
              else if (local_pf_num==0 && local_vf_num==1301 && local_vf_active==1) `fifo_error_check(1301)
              else if (local_pf_num==0 && local_vf_num==1302 && local_vf_active==1) `fifo_error_check(1302)
              else if (local_pf_num==0 && local_vf_num==1303 && local_vf_active==1) `fifo_error_check(1303)
              else if (local_pf_num==0 && local_vf_num==1304 && local_vf_active==1) `fifo_error_check(1304)
              else if (local_pf_num==0 && local_vf_num==1305 && local_vf_active==1) `fifo_error_check(1305)
              else if (local_pf_num==0 && local_vf_num==1306 && local_vf_active==1) `fifo_error_check(1306)
              else if (local_pf_num==0 && local_vf_num==1307 && local_vf_active==1) `fifo_error_check(1307)
              else if (local_pf_num==0 && local_vf_num==1308 && local_vf_active==1) `fifo_error_check(1308)
              else if (local_pf_num==0 && local_vf_num==1309 && local_vf_active==1) `fifo_error_check(1309)
              else if (local_pf_num==0 && local_vf_num==1310 && local_vf_active==1) `fifo_error_check(1310)
              else if (local_pf_num==0 && local_vf_num==1311 && local_vf_active==1) `fifo_error_check(1311)
              else if (local_pf_num==0 && local_vf_num==1312 && local_vf_active==1) `fifo_error_check(1312)
              else if (local_pf_num==0 && local_vf_num==1313 && local_vf_active==1) `fifo_error_check(1313)
              else if (local_pf_num==0 && local_vf_num==1314 && local_vf_active==1) `fifo_error_check(1314)
              else if (local_pf_num==0 && local_vf_num==1315 && local_vf_active==1) `fifo_error_check(1315)
              else if (local_pf_num==0 && local_vf_num==1316 && local_vf_active==1) `fifo_error_check(1316)
              else if (local_pf_num==0 && local_vf_num==1317 && local_vf_active==1) `fifo_error_check(1317)
              else if (local_pf_num==0 && local_vf_num==1318 && local_vf_active==1) `fifo_error_check(1318)
              else if (local_pf_num==0 && local_vf_num==1319 && local_vf_active==1) `fifo_error_check(1319)
              else if (local_pf_num==0 && local_vf_num==1320 && local_vf_active==1) `fifo_error_check(1320)
              else if (local_pf_num==0 && local_vf_num==1321 && local_vf_active==1) `fifo_error_check(1321)
              else if (local_pf_num==0 && local_vf_num==1322 && local_vf_active==1) `fifo_error_check(1322)
              else if (local_pf_num==0 && local_vf_num==1323 && local_vf_active==1) `fifo_error_check(1323)
              else if (local_pf_num==0 && local_vf_num==1324 && local_vf_active==1) `fifo_error_check(1324)
              else if (local_pf_num==0 && local_vf_num==1325 && local_vf_active==1) `fifo_error_check(1325)
              else if (local_pf_num==0 && local_vf_num==1326 && local_vf_active==1) `fifo_error_check(1326)
              else if (local_pf_num==0 && local_vf_num==1327 && local_vf_active==1) `fifo_error_check(1327)
              else if (local_pf_num==0 && local_vf_num==1328 && local_vf_active==1) `fifo_error_check(1328)
              else if (local_pf_num==0 && local_vf_num==1329 && local_vf_active==1) `fifo_error_check(1329)
              else if (local_pf_num==0 && local_vf_num==1330 && local_vf_active==1) `fifo_error_check(1330)
              else if (local_pf_num==0 && local_vf_num==1331 && local_vf_active==1) `fifo_error_check(1331)
              else if (local_pf_num==0 && local_vf_num==1332 && local_vf_active==1) `fifo_error_check(1332)
              else if (local_pf_num==0 && local_vf_num==1333 && local_vf_active==1) `fifo_error_check(1333)
              else if (local_pf_num==0 && local_vf_num==1334 && local_vf_active==1) `fifo_error_check(1334)
              else if (local_pf_num==0 && local_vf_num==1335 && local_vf_active==1) `fifo_error_check(1335)
              else if (local_pf_num==0 && local_vf_num==1336 && local_vf_active==1) `fifo_error_check(1336)
              else if (local_pf_num==0 && local_vf_num==1337 && local_vf_active==1) `fifo_error_check(1337)
              else if (local_pf_num==0 && local_vf_num==1338 && local_vf_active==1) `fifo_error_check(1338)
              else if (local_pf_num==0 && local_vf_num==1339 && local_vf_active==1) `fifo_error_check(1339)
              else if (local_pf_num==0 && local_vf_num==1340 && local_vf_active==1) `fifo_error_check(1340)
              else if (local_pf_num==0 && local_vf_num==1341 && local_vf_active==1) `fifo_error_check(1341)
              else if (local_pf_num==0 && local_vf_num==1342 && local_vf_active==1) `fifo_error_check(1342)
              else if (local_pf_num==0 && local_vf_num==1343 && local_vf_active==1) `fifo_error_check(1343)
              else if (local_pf_num==0 && local_vf_num==1344 && local_vf_active==1) `fifo_error_check(1344)
              else if (local_pf_num==0 && local_vf_num==1345 && local_vf_active==1) `fifo_error_check(1345)
              else if (local_pf_num==0 && local_vf_num==1346 && local_vf_active==1) `fifo_error_check(1346)
              else if (local_pf_num==0 && local_vf_num==1347 && local_vf_active==1) `fifo_error_check(1347)
              else if (local_pf_num==0 && local_vf_num==1348 && local_vf_active==1) `fifo_error_check(1348)
              else if (local_pf_num==0 && local_vf_num==1349 && local_vf_active==1) `fifo_error_check(1349)
              else if (local_pf_num==0 && local_vf_num==1350 && local_vf_active==1) `fifo_error_check(1350)
              else if (local_pf_num==0 && local_vf_num==1351 && local_vf_active==1) `fifo_error_check(1351)
              else if (local_pf_num==0 && local_vf_num==1352 && local_vf_active==1) `fifo_error_check(1352)
              else if (local_pf_num==0 && local_vf_num==1353 && local_vf_active==1) `fifo_error_check(1353)
              else if (local_pf_num==0 && local_vf_num==1354 && local_vf_active==1) `fifo_error_check(1354)
              else if (local_pf_num==0 && local_vf_num==1355 && local_vf_active==1) `fifo_error_check(1355)
              else if (local_pf_num==0 && local_vf_num==1356 && local_vf_active==1) `fifo_error_check(1356)
              else if (local_pf_num==0 && local_vf_num==1357 && local_vf_active==1) `fifo_error_check(1357)
              else if (local_pf_num==0 && local_vf_num==1358 && local_vf_active==1) `fifo_error_check(1358)
              else if (local_pf_num==0 && local_vf_num==1359 && local_vf_active==1) `fifo_error_check(1359)
              else if (local_pf_num==0 && local_vf_num==1360 && local_vf_active==1) `fifo_error_check(1360)
              else if (local_pf_num==0 && local_vf_num==1361 && local_vf_active==1) `fifo_error_check(1361)
              else if (local_pf_num==0 && local_vf_num==1362 && local_vf_active==1) `fifo_error_check(1362)
              else if (local_pf_num==0 && local_vf_num==1363 && local_vf_active==1) `fifo_error_check(1363)
              else if (local_pf_num==0 && local_vf_num==1364 && local_vf_active==1) `fifo_error_check(1364)
              else if (local_pf_num==0 && local_vf_num==1365 && local_vf_active==1) `fifo_error_check(1365)
              else if (local_pf_num==0 && local_vf_num==1366 && local_vf_active==1) `fifo_error_check(1366)
              else if (local_pf_num==0 && local_vf_num==1367 && local_vf_active==1) `fifo_error_check(1367)
              else if (local_pf_num==0 && local_vf_num==1368 && local_vf_active==1) `fifo_error_check(1368)
              else if (local_pf_num==0 && local_vf_num==1369 && local_vf_active==1) `fifo_error_check(1369)
              else if (local_pf_num==0 && local_vf_num==1370 && local_vf_active==1) `fifo_error_check(1370)
              else if (local_pf_num==0 && local_vf_num==1371 && local_vf_active==1) `fifo_error_check(1371)
              else if (local_pf_num==0 && local_vf_num==1372 && local_vf_active==1) `fifo_error_check(1372)
              else if (local_pf_num==0 && local_vf_num==1373 && local_vf_active==1) `fifo_error_check(1373)
              else if (local_pf_num==0 && local_vf_num==1374 && local_vf_active==1) `fifo_error_check(1374)
              else if (local_pf_num==0 && local_vf_num==1375 && local_vf_active==1) `fifo_error_check(1375)
              else if (local_pf_num==0 && local_vf_num==1376 && local_vf_active==1) `fifo_error_check(1376)
              else if (local_pf_num==0 && local_vf_num==1377 && local_vf_active==1) `fifo_error_check(1377)
              else if (local_pf_num==0 && local_vf_num==1378 && local_vf_active==1) `fifo_error_check(1378)
              else if (local_pf_num==0 && local_vf_num==1379 && local_vf_active==1) `fifo_error_check(1379)
              else if (local_pf_num==0 && local_vf_num==1380 && local_vf_active==1) `fifo_error_check(1380)
              else if (local_pf_num==0 && local_vf_num==1381 && local_vf_active==1) `fifo_error_check(1381)
              else if (local_pf_num==0 && local_vf_num==1382 && local_vf_active==1) `fifo_error_check(1382)
              else if (local_pf_num==0 && local_vf_num==1383 && local_vf_active==1) `fifo_error_check(1383)
              else if (local_pf_num==0 && local_vf_num==1384 && local_vf_active==1) `fifo_error_check(1384)
              else if (local_pf_num==0 && local_vf_num==1385 && local_vf_active==1) `fifo_error_check(1385)
              else if (local_pf_num==0 && local_vf_num==1386 && local_vf_active==1) `fifo_error_check(1386)
              else if (local_pf_num==0 && local_vf_num==1387 && local_vf_active==1) `fifo_error_check(1387)
              else if (local_pf_num==0 && local_vf_num==1388 && local_vf_active==1) `fifo_error_check(1388)
              else if (local_pf_num==0 && local_vf_num==1389 && local_vf_active==1) `fifo_error_check(1389)
              else if (local_pf_num==0 && local_vf_num==1390 && local_vf_active==1) `fifo_error_check(1390)
              else if (local_pf_num==0 && local_vf_num==1391 && local_vf_active==1) `fifo_error_check(1391)
              else if (local_pf_num==0 && local_vf_num==1392 && local_vf_active==1) `fifo_error_check(1392)
              else if (local_pf_num==0 && local_vf_num==1393 && local_vf_active==1) `fifo_error_check(1393)
              else if (local_pf_num==0 && local_vf_num==1394 && local_vf_active==1) `fifo_error_check(1394)
              else if (local_pf_num==0 && local_vf_num==1395 && local_vf_active==1) `fifo_error_check(1395)
              else if (local_pf_num==0 && local_vf_num==1396 && local_vf_active==1) `fifo_error_check(1396)
              else if (local_pf_num==0 && local_vf_num==1397 && local_vf_active==1) `fifo_error_check(1397)
              else if (local_pf_num==0 && local_vf_num==1398 && local_vf_active==1) `fifo_error_check(1398)
              else if (local_pf_num==0 && local_vf_num==1399 && local_vf_active==1) `fifo_error_check(1399)
              else if (local_pf_num==0 && local_vf_num==1400 && local_vf_active==1) `fifo_error_check(1400)
              else if (local_pf_num==0 && local_vf_num==1401 && local_vf_active==1) `fifo_error_check(1401)
              else if (local_pf_num==0 && local_vf_num==1402 && local_vf_active==1) `fifo_error_check(1402)
              else if (local_pf_num==0 && local_vf_num==1403 && local_vf_active==1) `fifo_error_check(1403)
              else if (local_pf_num==0 && local_vf_num==1404 && local_vf_active==1) `fifo_error_check(1404)
              else if (local_pf_num==0 && local_vf_num==1405 && local_vf_active==1) `fifo_error_check(1405)
              else if (local_pf_num==0 && local_vf_num==1406 && local_vf_active==1) `fifo_error_check(1406)
              else if (local_pf_num==0 && local_vf_num==1407 && local_vf_active==1) `fifo_error_check(1407)
              else if (local_pf_num==0 && local_vf_num==1408 && local_vf_active==1) `fifo_error_check(1408)
              else if (local_pf_num==0 && local_vf_num==1409 && local_vf_active==1) `fifo_error_check(1409)
              else if (local_pf_num==0 && local_vf_num==1410 && local_vf_active==1) `fifo_error_check(1410)
              else if (local_pf_num==0 && local_vf_num==1411 && local_vf_active==1) `fifo_error_check(1411)
              else if (local_pf_num==0 && local_vf_num==1412 && local_vf_active==1) `fifo_error_check(1412)
              else if (local_pf_num==0 && local_vf_num==1413 && local_vf_active==1) `fifo_error_check(1413)
              else if (local_pf_num==0 && local_vf_num==1414 && local_vf_active==1) `fifo_error_check(1414)
              else if (local_pf_num==0 && local_vf_num==1415 && local_vf_active==1) `fifo_error_check(1415)
              else if (local_pf_num==0 && local_vf_num==1416 && local_vf_active==1) `fifo_error_check(1416)
              else if (local_pf_num==0 && local_vf_num==1417 && local_vf_active==1) `fifo_error_check(1417)
              else if (local_pf_num==0 && local_vf_num==1418 && local_vf_active==1) `fifo_error_check(1418)
              else if (local_pf_num==0 && local_vf_num==1419 && local_vf_active==1) `fifo_error_check(1419)
              else if (local_pf_num==0 && local_vf_num==1420 && local_vf_active==1) `fifo_error_check(1420)
              else if (local_pf_num==0 && local_vf_num==1421 && local_vf_active==1) `fifo_error_check(1421)
              else if (local_pf_num==0 && local_vf_num==1422 && local_vf_active==1) `fifo_error_check(1422)
              else if (local_pf_num==0 && local_vf_num==1423 && local_vf_active==1) `fifo_error_check(1423)
              else if (local_pf_num==0 && local_vf_num==1424 && local_vf_active==1) `fifo_error_check(1424)
              else if (local_pf_num==0 && local_vf_num==1425 && local_vf_active==1) `fifo_error_check(1425)
              else if (local_pf_num==0 && local_vf_num==1426 && local_vf_active==1) `fifo_error_check(1426)
              else if (local_pf_num==0 && local_vf_num==1427 && local_vf_active==1) `fifo_error_check(1427)
              else if (local_pf_num==0 && local_vf_num==1428 && local_vf_active==1) `fifo_error_check(1428)
              else if (local_pf_num==0 && local_vf_num==1429 && local_vf_active==1) `fifo_error_check(1429)
              else if (local_pf_num==0 && local_vf_num==1430 && local_vf_active==1) `fifo_error_check(1430)
              else if (local_pf_num==0 && local_vf_num==1431 && local_vf_active==1) `fifo_error_check(1431)
              else if (local_pf_num==0 && local_vf_num==1432 && local_vf_active==1) `fifo_error_check(1432)
              else if (local_pf_num==0 && local_vf_num==1433 && local_vf_active==1) `fifo_error_check(1433)
              else if (local_pf_num==0 && local_vf_num==1434 && local_vf_active==1) `fifo_error_check(1434)
              else if (local_pf_num==0 && local_vf_num==1435 && local_vf_active==1) `fifo_error_check(1435)
              else if (local_pf_num==0 && local_vf_num==1436 && local_vf_active==1) `fifo_error_check(1436)
              else if (local_pf_num==0 && local_vf_num==1437 && local_vf_active==1) `fifo_error_check(1437)
              else if (local_pf_num==0 && local_vf_num==1438 && local_vf_active==1) `fifo_error_check(1438)
              else if (local_pf_num==0 && local_vf_num==1439 && local_vf_active==1) `fifo_error_check(1439)
              else if (local_pf_num==0 && local_vf_num==1440 && local_vf_active==1) `fifo_error_check(1440)
              else if (local_pf_num==0 && local_vf_num==1441 && local_vf_active==1) `fifo_error_check(1441)
              else if (local_pf_num==0 && local_vf_num==1442 && local_vf_active==1) `fifo_error_check(1442)
              else if (local_pf_num==0 && local_vf_num==1443 && local_vf_active==1) `fifo_error_check(1443)
              else if (local_pf_num==0 && local_vf_num==1444 && local_vf_active==1) `fifo_error_check(1444)
              else if (local_pf_num==0 && local_vf_num==1445 && local_vf_active==1) `fifo_error_check(1445)
              else if (local_pf_num==0 && local_vf_num==1446 && local_vf_active==1) `fifo_error_check(1446)
              else if (local_pf_num==0 && local_vf_num==1447 && local_vf_active==1) `fifo_error_check(1447)
              else if (local_pf_num==0 && local_vf_num==1448 && local_vf_active==1) `fifo_error_check(1448)
              else if (local_pf_num==0 && local_vf_num==1449 && local_vf_active==1) `fifo_error_check(1449)
              else if (local_pf_num==0 && local_vf_num==1450 && local_vf_active==1) `fifo_error_check(1450)
              else if (local_pf_num==0 && local_vf_num==1451 && local_vf_active==1) `fifo_error_check(1451)
              else if (local_pf_num==0 && local_vf_num==1452 && local_vf_active==1) `fifo_error_check(1452)
              else if (local_pf_num==0 && local_vf_num==1453 && local_vf_active==1) `fifo_error_check(1453)
              else if (local_pf_num==0 && local_vf_num==1454 && local_vf_active==1) `fifo_error_check(1454)
              else if (local_pf_num==0 && local_vf_num==1455 && local_vf_active==1) `fifo_error_check(1455)
              else if (local_pf_num==0 && local_vf_num==1456 && local_vf_active==1) `fifo_error_check(1456)
              else if (local_pf_num==0 && local_vf_num==1457 && local_vf_active==1) `fifo_error_check(1457)
              else if (local_pf_num==0 && local_vf_num==1458 && local_vf_active==1) `fifo_error_check(1458)
              else if (local_pf_num==0 && local_vf_num==1459 && local_vf_active==1) `fifo_error_check(1459)
              else if (local_pf_num==0 && local_vf_num==1460 && local_vf_active==1) `fifo_error_check(1460)
              else if (local_pf_num==0 && local_vf_num==1461 && local_vf_active==1) `fifo_error_check(1461)
              else if (local_pf_num==0 && local_vf_num==1462 && local_vf_active==1) `fifo_error_check(1462)
              else if (local_pf_num==0 && local_vf_num==1463 && local_vf_active==1) `fifo_error_check(1463)
              else if (local_pf_num==0 && local_vf_num==1464 && local_vf_active==1) `fifo_error_check(1464)
              else if (local_pf_num==0 && local_vf_num==1465 && local_vf_active==1) `fifo_error_check(1465)
              else if (local_pf_num==0 && local_vf_num==1466 && local_vf_active==1) `fifo_error_check(1466)
              else if (local_pf_num==0 && local_vf_num==1467 && local_vf_active==1) `fifo_error_check(1467)
              else if (local_pf_num==0 && local_vf_num==1468 && local_vf_active==1) `fifo_error_check(1468)
              else if (local_pf_num==0 && local_vf_num==1469 && local_vf_active==1) `fifo_error_check(1469)
              else if (local_pf_num==0 && local_vf_num==1470 && local_vf_active==1) `fifo_error_check(1470)
              else if (local_pf_num==0 && local_vf_num==1471 && local_vf_active==1) `fifo_error_check(1471)
              else if (local_pf_num==0 && local_vf_num==1472 && local_vf_active==1) `fifo_error_check(1472)
              else if (local_pf_num==0 && local_vf_num==1473 && local_vf_active==1) `fifo_error_check(1473)
              else if (local_pf_num==0 && local_vf_num==1474 && local_vf_active==1) `fifo_error_check(1474)
              else if (local_pf_num==0 && local_vf_num==1475 && local_vf_active==1) `fifo_error_check(1475)
              else if (local_pf_num==0 && local_vf_num==1476 && local_vf_active==1) `fifo_error_check(1476)
              else if (local_pf_num==0 && local_vf_num==1477 && local_vf_active==1) `fifo_error_check(1477)
              else if (local_pf_num==0 && local_vf_num==1478 && local_vf_active==1) `fifo_error_check(1478)
              else if (local_pf_num==0 && local_vf_num==1479 && local_vf_active==1) `fifo_error_check(1479)
              else if (local_pf_num==0 && local_vf_num==1480 && local_vf_active==1) `fifo_error_check(1480)
              else if (local_pf_num==0 && local_vf_num==1481 && local_vf_active==1) `fifo_error_check(1481)
              else if (local_pf_num==0 && local_vf_num==1482 && local_vf_active==1) `fifo_error_check(1482)
              else if (local_pf_num==0 && local_vf_num==1483 && local_vf_active==1) `fifo_error_check(1483)
              else if (local_pf_num==0 && local_vf_num==1484 && local_vf_active==1) `fifo_error_check(1484)
              else if (local_pf_num==0 && local_vf_num==1485 && local_vf_active==1) `fifo_error_check(1485)
              else if (local_pf_num==0 && local_vf_num==1486 && local_vf_active==1) `fifo_error_check(1486)
              else if (local_pf_num==0 && local_vf_num==1487 && local_vf_active==1) `fifo_error_check(1487)
              else if (local_pf_num==0 && local_vf_num==1488 && local_vf_active==1) `fifo_error_check(1488)
              else if (local_pf_num==0 && local_vf_num==1489 && local_vf_active==1) `fifo_error_check(1489)
              else if (local_pf_num==0 && local_vf_num==1490 && local_vf_active==1) `fifo_error_check(1490)
              else if (local_pf_num==0 && local_vf_num==1491 && local_vf_active==1) `fifo_error_check(1491)
              else if (local_pf_num==0 && local_vf_num==1492 && local_vf_active==1) `fifo_error_check(1492)
              else if (local_pf_num==0 && local_vf_num==1493 && local_vf_active==1) `fifo_error_check(1493)
              else if (local_pf_num==0 && local_vf_num==1494 && local_vf_active==1) `fifo_error_check(1494)
              else if (local_pf_num==0 && local_vf_num==1495 && local_vf_active==1) `fifo_error_check(1495)
              else if (local_pf_num==0 && local_vf_num==1496 && local_vf_active==1) `fifo_error_check(1496)
              else if (local_pf_num==0 && local_vf_num==1497 && local_vf_active==1) `fifo_error_check(1497)
              else if (local_pf_num==0 && local_vf_num==1498 && local_vf_active==1) `fifo_error_check(1498)
              else if (local_pf_num==0 && local_vf_num==1499 && local_vf_active==1) `fifo_error_check(1499)
              else if (local_pf_num==0 && local_vf_num==1500 && local_vf_active==1) `fifo_error_check(1500)
              else if (local_pf_num==0 && local_vf_num==1501 && local_vf_active==1) `fifo_error_check(1501)
              else if (local_pf_num==0 && local_vf_num==1502 && local_vf_active==1) `fifo_error_check(1502)
              else if (local_pf_num==0 && local_vf_num==1503 && local_vf_active==1) `fifo_error_check(1503)
              else if (local_pf_num==0 && local_vf_num==1504 && local_vf_active==1) `fifo_error_check(1504)
              else if (local_pf_num==0 && local_vf_num==1505 && local_vf_active==1) `fifo_error_check(1505)
              else if (local_pf_num==0 && local_vf_num==1506 && local_vf_active==1) `fifo_error_check(1506)
              else if (local_pf_num==0 && local_vf_num==1507 && local_vf_active==1) `fifo_error_check(1507)
              else if (local_pf_num==0 && local_vf_num==1508 && local_vf_active==1) `fifo_error_check(1508)
              else if (local_pf_num==0 && local_vf_num==1509 && local_vf_active==1) `fifo_error_check(1509)
              else if (local_pf_num==0 && local_vf_num==1510 && local_vf_active==1) `fifo_error_check(1510)
              else if (local_pf_num==0 && local_vf_num==1511 && local_vf_active==1) `fifo_error_check(1511)
              else if (local_pf_num==0 && local_vf_num==1512 && local_vf_active==1) `fifo_error_check(1512)
              else if (local_pf_num==0 && local_vf_num==1513 && local_vf_active==1) `fifo_error_check(1513)
              else if (local_pf_num==0 && local_vf_num==1514 && local_vf_active==1) `fifo_error_check(1514)
              else if (local_pf_num==0 && local_vf_num==1515 && local_vf_active==1) `fifo_error_check(1515)
              else if (local_pf_num==0 && local_vf_num==1516 && local_vf_active==1) `fifo_error_check(1516)
              else if (local_pf_num==0 && local_vf_num==1517 && local_vf_active==1) `fifo_error_check(1517)
              else if (local_pf_num==0 && local_vf_num==1518 && local_vf_active==1) `fifo_error_check(1518)
              else if (local_pf_num==0 && local_vf_num==1519 && local_vf_active==1) `fifo_error_check(1519)
              else if (local_pf_num==0 && local_vf_num==1520 && local_vf_active==1) `fifo_error_check(1520)
              else if (local_pf_num==0 && local_vf_num==1521 && local_vf_active==1) `fifo_error_check(1521)
              else if (local_pf_num==0 && local_vf_num==1522 && local_vf_active==1) `fifo_error_check(1522)
              else if (local_pf_num==0 && local_vf_num==1523 && local_vf_active==1) `fifo_error_check(1523)
              else if (local_pf_num==0 && local_vf_num==1524 && local_vf_active==1) `fifo_error_check(1524)
              else if (local_pf_num==0 && local_vf_num==1525 && local_vf_active==1) `fifo_error_check(1525)
              else if (local_pf_num==0 && local_vf_num==1526 && local_vf_active==1) `fifo_error_check(1526)
              else if (local_pf_num==0 && local_vf_num==1527 && local_vf_active==1) `fifo_error_check(1527)
              else if (local_pf_num==0 && local_vf_num==1528 && local_vf_active==1) `fifo_error_check(1528)
              else if (local_pf_num==0 && local_vf_num==1529 && local_vf_active==1) `fifo_error_check(1529)
              else if (local_pf_num==0 && local_vf_num==1530 && local_vf_active==1) `fifo_error_check(1530)
              else if (local_pf_num==0 && local_vf_num==1531 && local_vf_active==1) `fifo_error_check(1531)
              else if (local_pf_num==0 && local_vf_num==1532 && local_vf_active==1) `fifo_error_check(1532)
              else if (local_pf_num==0 && local_vf_num==1533 && local_vf_active==1) `fifo_error_check(1533)
              else if (local_pf_num==0 && local_vf_num==1534 && local_vf_active==1) `fifo_error_check(1534)
              else if (local_pf_num==0 && local_vf_num==1535 && local_vf_active==1) `fifo_error_check(1535)
              else if (local_pf_num==0 && local_vf_num==1536 && local_vf_active==1) `fifo_error_check(1536)
              else if (local_pf_num==0 && local_vf_num==1537 && local_vf_active==1) `fifo_error_check(1537)
              else if (local_pf_num==0 && local_vf_num==1538 && local_vf_active==1) `fifo_error_check(1538)
              else if (local_pf_num==0 && local_vf_num==1539 && local_vf_active==1) `fifo_error_check(1539)
              else if (local_pf_num==0 && local_vf_num==1540 && local_vf_active==1) `fifo_error_check(1540)
              else if (local_pf_num==0 && local_vf_num==1541 && local_vf_active==1) `fifo_error_check(1541)
              else if (local_pf_num==0 && local_vf_num==1542 && local_vf_active==1) `fifo_error_check(1542)
              else if (local_pf_num==0 && local_vf_num==1543 && local_vf_active==1) `fifo_error_check(1543)
              else if (local_pf_num==0 && local_vf_num==1544 && local_vf_active==1) `fifo_error_check(1544)
              else if (local_pf_num==0 && local_vf_num==1545 && local_vf_active==1) `fifo_error_check(1545)
              else if (local_pf_num==0 && local_vf_num==1546 && local_vf_active==1) `fifo_error_check(1546)
              else if (local_pf_num==0 && local_vf_num==1547 && local_vf_active==1) `fifo_error_check(1547)
              else if (local_pf_num==0 && local_vf_num==1548 && local_vf_active==1) `fifo_error_check(1548)
              else if (local_pf_num==0 && local_vf_num==1549 && local_vf_active==1) `fifo_error_check(1549)
              else if (local_pf_num==0 && local_vf_num==1550 && local_vf_active==1) `fifo_error_check(1550)
              else if (local_pf_num==0 && local_vf_num==1551 && local_vf_active==1) `fifo_error_check(1551)
              else if (local_pf_num==0 && local_vf_num==1552 && local_vf_active==1) `fifo_error_check(1552)
              else if (local_pf_num==0 && local_vf_num==1553 && local_vf_active==1) `fifo_error_check(1553)
              else if (local_pf_num==0 && local_vf_num==1554 && local_vf_active==1) `fifo_error_check(1554)
              else if (local_pf_num==0 && local_vf_num==1555 && local_vf_active==1) `fifo_error_check(1555)
              else if (local_pf_num==0 && local_vf_num==1556 && local_vf_active==1) `fifo_error_check(1556)
              else if (local_pf_num==0 && local_vf_num==1557 && local_vf_active==1) `fifo_error_check(1557)
              else if (local_pf_num==0 && local_vf_num==1558 && local_vf_active==1) `fifo_error_check(1558)
              else if (local_pf_num==0 && local_vf_num==1559 && local_vf_active==1) `fifo_error_check(1559)
              else if (local_pf_num==0 && local_vf_num==1560 && local_vf_active==1) `fifo_error_check(1560)
              else if (local_pf_num==0 && local_vf_num==1561 && local_vf_active==1) `fifo_error_check(1561)
              else if (local_pf_num==0 && local_vf_num==1562 && local_vf_active==1) `fifo_error_check(1562)
              else if (local_pf_num==0 && local_vf_num==1563 && local_vf_active==1) `fifo_error_check(1563)
              else if (local_pf_num==0 && local_vf_num==1564 && local_vf_active==1) `fifo_error_check(1564)
              else if (local_pf_num==0 && local_vf_num==1565 && local_vf_active==1) `fifo_error_check(1565)
              else if (local_pf_num==0 && local_vf_num==1566 && local_vf_active==1) `fifo_error_check(1566)
              else if (local_pf_num==0 && local_vf_num==1567 && local_vf_active==1) `fifo_error_check(1567)
              else if (local_pf_num==0 && local_vf_num==1568 && local_vf_active==1) `fifo_error_check(1568)
              else if (local_pf_num==0 && local_vf_num==1569 && local_vf_active==1) `fifo_error_check(1569)
              else if (local_pf_num==0 && local_vf_num==1570 && local_vf_active==1) `fifo_error_check(1570)
              else if (local_pf_num==0 && local_vf_num==1571 && local_vf_active==1) `fifo_error_check(1571)
              else if (local_pf_num==0 && local_vf_num==1572 && local_vf_active==1) `fifo_error_check(1572)
              else if (local_pf_num==0 && local_vf_num==1573 && local_vf_active==1) `fifo_error_check(1573)
              else if (local_pf_num==0 && local_vf_num==1574 && local_vf_active==1) `fifo_error_check(1574)
              else if (local_pf_num==0 && local_vf_num==1575 && local_vf_active==1) `fifo_error_check(1575)
              else if (local_pf_num==0 && local_vf_num==1576 && local_vf_active==1) `fifo_error_check(1576)
              else if (local_pf_num==0 && local_vf_num==1577 && local_vf_active==1) `fifo_error_check(1577)
              else if (local_pf_num==0 && local_vf_num==1578 && local_vf_active==1) `fifo_error_check(1578)
              else if (local_pf_num==0 && local_vf_num==1579 && local_vf_active==1) `fifo_error_check(1579)
              else if (local_pf_num==0 && local_vf_num==1580 && local_vf_active==1) `fifo_error_check(1580)
              else if (local_pf_num==0 && local_vf_num==1581 && local_vf_active==1) `fifo_error_check(1581)
              else if (local_pf_num==0 && local_vf_num==1582 && local_vf_active==1) `fifo_error_check(1582)
              else if (local_pf_num==0 && local_vf_num==1583 && local_vf_active==1) `fifo_error_check(1583)
              else if (local_pf_num==0 && local_vf_num==1584 && local_vf_active==1) `fifo_error_check(1584)
              else if (local_pf_num==0 && local_vf_num==1585 && local_vf_active==1) `fifo_error_check(1585)
              else if (local_pf_num==0 && local_vf_num==1586 && local_vf_active==1) `fifo_error_check(1586)
              else if (local_pf_num==0 && local_vf_num==1587 && local_vf_active==1) `fifo_error_check(1587)
              else if (local_pf_num==0 && local_vf_num==1588 && local_vf_active==1) `fifo_error_check(1588)
              else if (local_pf_num==0 && local_vf_num==1589 && local_vf_active==1) `fifo_error_check(1589)
              else if (local_pf_num==0 && local_vf_num==1590 && local_vf_active==1) `fifo_error_check(1590)
              else if (local_pf_num==0 && local_vf_num==1591 && local_vf_active==1) `fifo_error_check(1591)
              else if (local_pf_num==0 && local_vf_num==1592 && local_vf_active==1) `fifo_error_check(1592)
              else if (local_pf_num==0 && local_vf_num==1593 && local_vf_active==1) `fifo_error_check(1593)
              else if (local_pf_num==0 && local_vf_num==1594 && local_vf_active==1) `fifo_error_check(1594)
              else if (local_pf_num==0 && local_vf_num==1595 && local_vf_active==1) `fifo_error_check(1595)
              else if (local_pf_num==0 && local_vf_num==1596 && local_vf_active==1) `fifo_error_check(1596)
              else if (local_pf_num==0 && local_vf_num==1597 && local_vf_active==1) `fifo_error_check(1597)
              else if (local_pf_num==0 && local_vf_num==1598 && local_vf_active==1) `fifo_error_check(1598)
              else if (local_pf_num==0 && local_vf_num==1599 && local_vf_active==1) `fifo_error_check(1599)
              else if (local_pf_num==0 && local_vf_num==1600 && local_vf_active==1) `fifo_error_check(1600)
              else if (local_pf_num==0 && local_vf_num==1601 && local_vf_active==1) `fifo_error_check(1601)
              else if (local_pf_num==0 && local_vf_num==1602 && local_vf_active==1) `fifo_error_check(1602)
              else if (local_pf_num==0 && local_vf_num==1603 && local_vf_active==1) `fifo_error_check(1603)
              else if (local_pf_num==0 && local_vf_num==1604 && local_vf_active==1) `fifo_error_check(1604)
              else if (local_pf_num==0 && local_vf_num==1605 && local_vf_active==1) `fifo_error_check(1605)
              else if (local_pf_num==0 && local_vf_num==1606 && local_vf_active==1) `fifo_error_check(1606)
              else if (local_pf_num==0 && local_vf_num==1607 && local_vf_active==1) `fifo_error_check(1607)
              else if (local_pf_num==0 && local_vf_num==1608 && local_vf_active==1) `fifo_error_check(1608)
              else if (local_pf_num==0 && local_vf_num==1609 && local_vf_active==1) `fifo_error_check(1609)
              else if (local_pf_num==0 && local_vf_num==1610 && local_vf_active==1) `fifo_error_check(1610)
              else if (local_pf_num==0 && local_vf_num==1611 && local_vf_active==1) `fifo_error_check(1611)
              else if (local_pf_num==0 && local_vf_num==1612 && local_vf_active==1) `fifo_error_check(1612)
              else if (local_pf_num==0 && local_vf_num==1613 && local_vf_active==1) `fifo_error_check(1613)
              else if (local_pf_num==0 && local_vf_num==1614 && local_vf_active==1) `fifo_error_check(1614)
              else if (local_pf_num==0 && local_vf_num==1615 && local_vf_active==1) `fifo_error_check(1615)
              else if (local_pf_num==0 && local_vf_num==1616 && local_vf_active==1) `fifo_error_check(1616)
              else if (local_pf_num==0 && local_vf_num==1617 && local_vf_active==1) `fifo_error_check(1617)
              else if (local_pf_num==0 && local_vf_num==1618 && local_vf_active==1) `fifo_error_check(1618)
              else if (local_pf_num==0 && local_vf_num==1619 && local_vf_active==1) `fifo_error_check(1619)
              else if (local_pf_num==0 && local_vf_num==1620 && local_vf_active==1) `fifo_error_check(1620)
              else if (local_pf_num==0 && local_vf_num==1621 && local_vf_active==1) `fifo_error_check(1621)
              else if (local_pf_num==0 && local_vf_num==1622 && local_vf_active==1) `fifo_error_check(1622)
              else if (local_pf_num==0 && local_vf_num==1623 && local_vf_active==1) `fifo_error_check(1623)
              else if (local_pf_num==0 && local_vf_num==1624 && local_vf_active==1) `fifo_error_check(1624)
              else if (local_pf_num==0 && local_vf_num==1625 && local_vf_active==1) `fifo_error_check(1625)
              else if (local_pf_num==0 && local_vf_num==1626 && local_vf_active==1) `fifo_error_check(1626)
              else if (local_pf_num==0 && local_vf_num==1627 && local_vf_active==1) `fifo_error_check(1627)
              else if (local_pf_num==0 && local_vf_num==1628 && local_vf_active==1) `fifo_error_check(1628)
              else if (local_pf_num==0 && local_vf_num==1629 && local_vf_active==1) `fifo_error_check(1629)
              else if (local_pf_num==0 && local_vf_num==1630 && local_vf_active==1) `fifo_error_check(1630)
              else if (local_pf_num==0 && local_vf_num==1631 && local_vf_active==1) `fifo_error_check(1631)
              else if (local_pf_num==0 && local_vf_num==1632 && local_vf_active==1) `fifo_error_check(1632)
              else if (local_pf_num==0 && local_vf_num==1633 && local_vf_active==1) `fifo_error_check(1633)
              else if (local_pf_num==0 && local_vf_num==1634 && local_vf_active==1) `fifo_error_check(1634)
              else if (local_pf_num==0 && local_vf_num==1635 && local_vf_active==1) `fifo_error_check(1635)
              else if (local_pf_num==0 && local_vf_num==1636 && local_vf_active==1) `fifo_error_check(1636)
              else if (local_pf_num==0 && local_vf_num==1637 && local_vf_active==1) `fifo_error_check(1637)
              else if (local_pf_num==0 && local_vf_num==1638 && local_vf_active==1) `fifo_error_check(1638)
              else if (local_pf_num==0 && local_vf_num==1639 && local_vf_active==1) `fifo_error_check(1639)
              else if (local_pf_num==0 && local_vf_num==1640 && local_vf_active==1) `fifo_error_check(1640)
              else if (local_pf_num==0 && local_vf_num==1641 && local_vf_active==1) `fifo_error_check(1641)
              else if (local_pf_num==0 && local_vf_num==1642 && local_vf_active==1) `fifo_error_check(1642)
              else if (local_pf_num==0 && local_vf_num==1643 && local_vf_active==1) `fifo_error_check(1643)
              else if (local_pf_num==0 && local_vf_num==1644 && local_vf_active==1) `fifo_error_check(1644)
              else if (local_pf_num==0 && local_vf_num==1645 && local_vf_active==1) `fifo_error_check(1645)
              else if (local_pf_num==0 && local_vf_num==1646 && local_vf_active==1) `fifo_error_check(1646)
              else if (local_pf_num==0 && local_vf_num==1647 && local_vf_active==1) `fifo_error_check(1647)
              else if (local_pf_num==0 && local_vf_num==1648 && local_vf_active==1) `fifo_error_check(1648)
              else if (local_pf_num==0 && local_vf_num==1649 && local_vf_active==1) `fifo_error_check(1649)
              else if (local_pf_num==0 && local_vf_num==1650 && local_vf_active==1) `fifo_error_check(1650)
              else if (local_pf_num==0 && local_vf_num==1651 && local_vf_active==1) `fifo_error_check(1651)
              else if (local_pf_num==0 && local_vf_num==1652 && local_vf_active==1) `fifo_error_check(1652)
              else if (local_pf_num==0 && local_vf_num==1653 && local_vf_active==1) `fifo_error_check(1653)
              else if (local_pf_num==0 && local_vf_num==1654 && local_vf_active==1) `fifo_error_check(1654)
              else if (local_pf_num==0 && local_vf_num==1655 && local_vf_active==1) `fifo_error_check(1655)
              else if (local_pf_num==0 && local_vf_num==1656 && local_vf_active==1) `fifo_error_check(1656)
              else if (local_pf_num==0 && local_vf_num==1657 && local_vf_active==1) `fifo_error_check(1657)
              else if (local_pf_num==0 && local_vf_num==1658 && local_vf_active==1) `fifo_error_check(1658)
              else if (local_pf_num==0 && local_vf_num==1659 && local_vf_active==1) `fifo_error_check(1659)
              else if (local_pf_num==0 && local_vf_num==1660 && local_vf_active==1) `fifo_error_check(1660)
              else if (local_pf_num==0 && local_vf_num==1661 && local_vf_active==1) `fifo_error_check(1661)
              else if (local_pf_num==0 && local_vf_num==1662 && local_vf_active==1) `fifo_error_check(1662)
              else if (local_pf_num==0 && local_vf_num==1663 && local_vf_active==1) `fifo_error_check(1663)
              else if (local_pf_num==0 && local_vf_num==1664 && local_vf_active==1) `fifo_error_check(1664)
              else if (local_pf_num==0 && local_vf_num==1665 && local_vf_active==1) `fifo_error_check(1665)
              else if (local_pf_num==0 && local_vf_num==1666 && local_vf_active==1) `fifo_error_check(1666)
              else if (local_pf_num==0 && local_vf_num==1667 && local_vf_active==1) `fifo_error_check(1667)
              else if (local_pf_num==0 && local_vf_num==1668 && local_vf_active==1) `fifo_error_check(1668)
              else if (local_pf_num==0 && local_vf_num==1669 && local_vf_active==1) `fifo_error_check(1669)
              else if (local_pf_num==0 && local_vf_num==1670 && local_vf_active==1) `fifo_error_check(1670)
              else if (local_pf_num==0 && local_vf_num==1671 && local_vf_active==1) `fifo_error_check(1671)
              else if (local_pf_num==0 && local_vf_num==1672 && local_vf_active==1) `fifo_error_check(1672)
              else if (local_pf_num==0 && local_vf_num==1673 && local_vf_active==1) `fifo_error_check(1673)
              else if (local_pf_num==0 && local_vf_num==1674 && local_vf_active==1) `fifo_error_check(1674)
              else if (local_pf_num==0 && local_vf_num==1675 && local_vf_active==1) `fifo_error_check(1675)
              else if (local_pf_num==0 && local_vf_num==1676 && local_vf_active==1) `fifo_error_check(1676)
              else if (local_pf_num==0 && local_vf_num==1677 && local_vf_active==1) `fifo_error_check(1677)
              else if (local_pf_num==0 && local_vf_num==1678 && local_vf_active==1) `fifo_error_check(1678)
              else if (local_pf_num==0 && local_vf_num==1679 && local_vf_active==1) `fifo_error_check(1679)
              else if (local_pf_num==0 && local_vf_num==1680 && local_vf_active==1) `fifo_error_check(1680)
              else if (local_pf_num==0 && local_vf_num==1681 && local_vf_active==1) `fifo_error_check(1681)
              else if (local_pf_num==0 && local_vf_num==1682 && local_vf_active==1) `fifo_error_check(1682)
              else if (local_pf_num==0 && local_vf_num==1683 && local_vf_active==1) `fifo_error_check(1683)
              else if (local_pf_num==0 && local_vf_num==1684 && local_vf_active==1) `fifo_error_check(1684)
              else if (local_pf_num==0 && local_vf_num==1685 && local_vf_active==1) `fifo_error_check(1685)
              else if (local_pf_num==0 && local_vf_num==1686 && local_vf_active==1) `fifo_error_check(1686)
              else if (local_pf_num==0 && local_vf_num==1687 && local_vf_active==1) `fifo_error_check(1687)
              else if (local_pf_num==0 && local_vf_num==1688 && local_vf_active==1) `fifo_error_check(1688)
              else if (local_pf_num==0 && local_vf_num==1689 && local_vf_active==1) `fifo_error_check(1689)
              else if (local_pf_num==0 && local_vf_num==1690 && local_vf_active==1) `fifo_error_check(1690)
              else if (local_pf_num==0 && local_vf_num==1691 && local_vf_active==1) `fifo_error_check(1691)
              else if (local_pf_num==0 && local_vf_num==1692 && local_vf_active==1) `fifo_error_check(1692)
              else if (local_pf_num==0 && local_vf_num==1693 && local_vf_active==1) `fifo_error_check(1693)
              else if (local_pf_num==0 && local_vf_num==1694 && local_vf_active==1) `fifo_error_check(1694)
              else if (local_pf_num==0 && local_vf_num==1695 && local_vf_active==1) `fifo_error_check(1695)
              else if (local_pf_num==0 && local_vf_num==1696 && local_vf_active==1) `fifo_error_check(1696)
              else if (local_pf_num==0 && local_vf_num==1697 && local_vf_active==1) `fifo_error_check(1697)
              else if (local_pf_num==0 && local_vf_num==1698 && local_vf_active==1) `fifo_error_check(1698)
              else if (local_pf_num==0 && local_vf_num==1699 && local_vf_active==1) `fifo_error_check(1699)
              else if (local_pf_num==0 && local_vf_num==1700 && local_vf_active==1) `fifo_error_check(1700)
              else if (local_pf_num==0 && local_vf_num==1701 && local_vf_active==1) `fifo_error_check(1701)
              else if (local_pf_num==0 && local_vf_num==1702 && local_vf_active==1) `fifo_error_check(1702)
              else if (local_pf_num==0 && local_vf_num==1703 && local_vf_active==1) `fifo_error_check(1703)
              else if (local_pf_num==0 && local_vf_num==1704 && local_vf_active==1) `fifo_error_check(1704)
              else if (local_pf_num==0 && local_vf_num==1705 && local_vf_active==1) `fifo_error_check(1705)
              else if (local_pf_num==0 && local_vf_num==1706 && local_vf_active==1) `fifo_error_check(1706)
              else if (local_pf_num==0 && local_vf_num==1707 && local_vf_active==1) `fifo_error_check(1707)
              else if (local_pf_num==0 && local_vf_num==1708 && local_vf_active==1) `fifo_error_check(1708)
              else if (local_pf_num==0 && local_vf_num==1709 && local_vf_active==1) `fifo_error_check(1709)
              else if (local_pf_num==0 && local_vf_num==1710 && local_vf_active==1) `fifo_error_check(1710)
              else if (local_pf_num==0 && local_vf_num==1711 && local_vf_active==1) `fifo_error_check(1711)
              else if (local_pf_num==0 && local_vf_num==1712 && local_vf_active==1) `fifo_error_check(1712)
              else if (local_pf_num==0 && local_vf_num==1713 && local_vf_active==1) `fifo_error_check(1713)
              else if (local_pf_num==0 && local_vf_num==1714 && local_vf_active==1) `fifo_error_check(1714)
              else if (local_pf_num==0 && local_vf_num==1715 && local_vf_active==1) `fifo_error_check(1715)
              else if (local_pf_num==0 && local_vf_num==1716 && local_vf_active==1) `fifo_error_check(1716)
              else if (local_pf_num==0 && local_vf_num==1717 && local_vf_active==1) `fifo_error_check(1717)
              else if (local_pf_num==0 && local_vf_num==1718 && local_vf_active==1) `fifo_error_check(1718)
              else if (local_pf_num==0 && local_vf_num==1719 && local_vf_active==1) `fifo_error_check(1719)
              else if (local_pf_num==0 && local_vf_num==1720 && local_vf_active==1) `fifo_error_check(1720)
              else if (local_pf_num==0 && local_vf_num==1721 && local_vf_active==1) `fifo_error_check(1721)
              else if (local_pf_num==0 && local_vf_num==1722 && local_vf_active==1) `fifo_error_check(1722)
              else if (local_pf_num==0 && local_vf_num==1723 && local_vf_active==1) `fifo_error_check(1723)
              else if (local_pf_num==0 && local_vf_num==1724 && local_vf_active==1) `fifo_error_check(1724)
              else if (local_pf_num==0 && local_vf_num==1725 && local_vf_active==1) `fifo_error_check(1725)
              else if (local_pf_num==0 && local_vf_num==1726 && local_vf_active==1) `fifo_error_check(1726)
              else if (local_pf_num==0 && local_vf_num==1727 && local_vf_active==1) `fifo_error_check(1727)
              else if (local_pf_num==0 && local_vf_num==1728 && local_vf_active==1) `fifo_error_check(1728)
              else if (local_pf_num==0 && local_vf_num==1729 && local_vf_active==1) `fifo_error_check(1729)
              else if (local_pf_num==0 && local_vf_num==1730 && local_vf_active==1) `fifo_error_check(1730)
              else if (local_pf_num==0 && local_vf_num==1731 && local_vf_active==1) `fifo_error_check(1731)
              else if (local_pf_num==0 && local_vf_num==1732 && local_vf_active==1) `fifo_error_check(1732)
              else if (local_pf_num==0 && local_vf_num==1733 && local_vf_active==1) `fifo_error_check(1733)
              else if (local_pf_num==0 && local_vf_num==1734 && local_vf_active==1) `fifo_error_check(1734)
              else if (local_pf_num==0 && local_vf_num==1735 && local_vf_active==1) `fifo_error_check(1735)
              else if (local_pf_num==0 && local_vf_num==1736 && local_vf_active==1) `fifo_error_check(1736)
              else if (local_pf_num==0 && local_vf_num==1737 && local_vf_active==1) `fifo_error_check(1737)
              else if (local_pf_num==0 && local_vf_num==1738 && local_vf_active==1) `fifo_error_check(1738)
              else if (local_pf_num==0 && local_vf_num==1739 && local_vf_active==1) `fifo_error_check(1739)
              else if (local_pf_num==0 && local_vf_num==1740 && local_vf_active==1) `fifo_error_check(1740)
              else if (local_pf_num==0 && local_vf_num==1741 && local_vf_active==1) `fifo_error_check(1741)
              else if (local_pf_num==0 && local_vf_num==1742 && local_vf_active==1) `fifo_error_check(1742)
              else if (local_pf_num==0 && local_vf_num==1743 && local_vf_active==1) `fifo_error_check(1743)
              else if (local_pf_num==0 && local_vf_num==1744 && local_vf_active==1) `fifo_error_check(1744)
              else if (local_pf_num==0 && local_vf_num==1745 && local_vf_active==1) `fifo_error_check(1745)
              else if (local_pf_num==0 && local_vf_num==1746 && local_vf_active==1) `fifo_error_check(1746)
              else if (local_pf_num==0 && local_vf_num==1747 && local_vf_active==1) `fifo_error_check(1747)
              else if (local_pf_num==0 && local_vf_num==1748 && local_vf_active==1) `fifo_error_check(1748)
              else if (local_pf_num==0 && local_vf_num==1749 && local_vf_active==1) `fifo_error_check(1749)
              else if (local_pf_num==0 && local_vf_num==1750 && local_vf_active==1) `fifo_error_check(1750)
              else if (local_pf_num==0 && local_vf_num==1751 && local_vf_active==1) `fifo_error_check(1751)
              else if (local_pf_num==0 && local_vf_num==1752 && local_vf_active==1) `fifo_error_check(1752)
              else if (local_pf_num==0 && local_vf_num==1753 && local_vf_active==1) `fifo_error_check(1753)
              else if (local_pf_num==0 && local_vf_num==1754 && local_vf_active==1) `fifo_error_check(1754)
              else if (local_pf_num==0 && local_vf_num==1755 && local_vf_active==1) `fifo_error_check(1755)
              else if (local_pf_num==0 && local_vf_num==1756 && local_vf_active==1) `fifo_error_check(1756)
              else if (local_pf_num==0 && local_vf_num==1757 && local_vf_active==1) `fifo_error_check(1757)
              else if (local_pf_num==0 && local_vf_num==1758 && local_vf_active==1) `fifo_error_check(1758)
              else if (local_pf_num==0 && local_vf_num==1759 && local_vf_active==1) `fifo_error_check(1759)
              else if (local_pf_num==0 && local_vf_num==1760 && local_vf_active==1) `fifo_error_check(1760)
              else if (local_pf_num==0 && local_vf_num==1761 && local_vf_active==1) `fifo_error_check(1761)
              else if (local_pf_num==0 && local_vf_num==1762 && local_vf_active==1) `fifo_error_check(1762)
              else if (local_pf_num==0 && local_vf_num==1763 && local_vf_active==1) `fifo_error_check(1763)
              else if (local_pf_num==0 && local_vf_num==1764 && local_vf_active==1) `fifo_error_check(1764)
              else if (local_pf_num==0 && local_vf_num==1765 && local_vf_active==1) `fifo_error_check(1765)
              else if (local_pf_num==0 && local_vf_num==1766 && local_vf_active==1) `fifo_error_check(1766)
              else if (local_pf_num==0 && local_vf_num==1767 && local_vf_active==1) `fifo_error_check(1767)
              else if (local_pf_num==0 && local_vf_num==1768 && local_vf_active==1) `fifo_error_check(1768)
              else if (local_pf_num==0 && local_vf_num==1769 && local_vf_active==1) `fifo_error_check(1769)
              else if (local_pf_num==0 && local_vf_num==1770 && local_vf_active==1) `fifo_error_check(1770)
              else if (local_pf_num==0 && local_vf_num==1771 && local_vf_active==1) `fifo_error_check(1771)
              else if (local_pf_num==0 && local_vf_num==1772 && local_vf_active==1) `fifo_error_check(1772)
              else if (local_pf_num==0 && local_vf_num==1773 && local_vf_active==1) `fifo_error_check(1773)
              else if (local_pf_num==0 && local_vf_num==1774 && local_vf_active==1) `fifo_error_check(1774)
              else if (local_pf_num==0 && local_vf_num==1775 && local_vf_active==1) `fifo_error_check(1775)
              else if (local_pf_num==0 && local_vf_num==1776 && local_vf_active==1) `fifo_error_check(1776)
              else if (local_pf_num==0 && local_vf_num==1777 && local_vf_active==1) `fifo_error_check(1777)
              else if (local_pf_num==0 && local_vf_num==1778 && local_vf_active==1) `fifo_error_check(1778)
              else if (local_pf_num==0 && local_vf_num==1779 && local_vf_active==1) `fifo_error_check(1779)
              else if (local_pf_num==0 && local_vf_num==1780 && local_vf_active==1) `fifo_error_check(1780)
              else if (local_pf_num==0 && local_vf_num==1781 && local_vf_active==1) `fifo_error_check(1781)
              else if (local_pf_num==0 && local_vf_num==1782 && local_vf_active==1) `fifo_error_check(1782)
              else if (local_pf_num==0 && local_vf_num==1783 && local_vf_active==1) `fifo_error_check(1783)
              else if (local_pf_num==0 && local_vf_num==1784 && local_vf_active==1) `fifo_error_check(1784)
              else if (local_pf_num==0 && local_vf_num==1785 && local_vf_active==1) `fifo_error_check(1785)
              else if (local_pf_num==0 && local_vf_num==1786 && local_vf_active==1) `fifo_error_check(1786)
              else if (local_pf_num==0 && local_vf_num==1787 && local_vf_active==1) `fifo_error_check(1787)
              else if (local_pf_num==0 && local_vf_num==1788 && local_vf_active==1) `fifo_error_check(1788)
              else if (local_pf_num==0 && local_vf_num==1789 && local_vf_active==1) `fifo_error_check(1789)
              else if (local_pf_num==0 && local_vf_num==1790 && local_vf_active==1) `fifo_error_check(1790)
              else if (local_pf_num==0 && local_vf_num==1791 && local_vf_active==1) `fifo_error_check(1791)
              else if (local_pf_num==0 && local_vf_num==1792 && local_vf_active==1) `fifo_error_check(1792)
              else if (local_pf_num==0 && local_vf_num==1793 && local_vf_active==1) `fifo_error_check(1793)
              else if (local_pf_num==0 && local_vf_num==1794 && local_vf_active==1) `fifo_error_check(1794)
              else if (local_pf_num==0 && local_vf_num==1795 && local_vf_active==1) `fifo_error_check(1795)
              else if (local_pf_num==0 && local_vf_num==1796 && local_vf_active==1) `fifo_error_check(1796)
              else if (local_pf_num==0 && local_vf_num==1797 && local_vf_active==1) `fifo_error_check(1797)
              else if (local_pf_num==0 && local_vf_num==1798 && local_vf_active==1) `fifo_error_check(1798)
              else if (local_pf_num==0 && local_vf_num==1799 && local_vf_active==1) `fifo_error_check(1799)
              else if (local_pf_num==0 && local_vf_num==1800 && local_vf_active==1) `fifo_error_check(1800)
              else if (local_pf_num==0 && local_vf_num==1801 && local_vf_active==1) `fifo_error_check(1801)
              else if (local_pf_num==0 && local_vf_num==1802 && local_vf_active==1) `fifo_error_check(1802)
              else if (local_pf_num==0 && local_vf_num==1803 && local_vf_active==1) `fifo_error_check(1803)
              else if (local_pf_num==0 && local_vf_num==1804 && local_vf_active==1) `fifo_error_check(1804)
              else if (local_pf_num==0 && local_vf_num==1805 && local_vf_active==1) `fifo_error_check(1805)
              else if (local_pf_num==0 && local_vf_num==1806 && local_vf_active==1) `fifo_error_check(1806)
              else if (local_pf_num==0 && local_vf_num==1807 && local_vf_active==1) `fifo_error_check(1807)
              else if (local_pf_num==0 && local_vf_num==1808 && local_vf_active==1) `fifo_error_check(1808)
              else if (local_pf_num==0 && local_vf_num==1809 && local_vf_active==1) `fifo_error_check(1809)
              else if (local_pf_num==0 && local_vf_num==1810 && local_vf_active==1) `fifo_error_check(1810)
              else if (local_pf_num==0 && local_vf_num==1811 && local_vf_active==1) `fifo_error_check(1811)
              else if (local_pf_num==0 && local_vf_num==1812 && local_vf_active==1) `fifo_error_check(1812)
              else if (local_pf_num==0 && local_vf_num==1813 && local_vf_active==1) `fifo_error_check(1813)
              else if (local_pf_num==0 && local_vf_num==1814 && local_vf_active==1) `fifo_error_check(1814)
              else if (local_pf_num==0 && local_vf_num==1815 && local_vf_active==1) `fifo_error_check(1815)
              else if (local_pf_num==0 && local_vf_num==1816 && local_vf_active==1) `fifo_error_check(1816)
              else if (local_pf_num==0 && local_vf_num==1817 && local_vf_active==1) `fifo_error_check(1817)
              else if (local_pf_num==0 && local_vf_num==1818 && local_vf_active==1) `fifo_error_check(1818)
              else if (local_pf_num==0 && local_vf_num==1819 && local_vf_active==1) `fifo_error_check(1819)
              else if (local_pf_num==0 && local_vf_num==1820 && local_vf_active==1) `fifo_error_check(1820)
              else if (local_pf_num==0 && local_vf_num==1821 && local_vf_active==1) `fifo_error_check(1821)
              else if (local_pf_num==0 && local_vf_num==1822 && local_vf_active==1) `fifo_error_check(1822)
              else if (local_pf_num==0 && local_vf_num==1823 && local_vf_active==1) `fifo_error_check(1823)
              else if (local_pf_num==0 && local_vf_num==1824 && local_vf_active==1) `fifo_error_check(1824)
              else if (local_pf_num==0 && local_vf_num==1825 && local_vf_active==1) `fifo_error_check(1825)
              else if (local_pf_num==0 && local_vf_num==1826 && local_vf_active==1) `fifo_error_check(1826)
              else if (local_pf_num==0 && local_vf_num==1827 && local_vf_active==1) `fifo_error_check(1827)
              else if (local_pf_num==0 && local_vf_num==1828 && local_vf_active==1) `fifo_error_check(1828)
              else if (local_pf_num==0 && local_vf_num==1829 && local_vf_active==1) `fifo_error_check(1829)
              else if (local_pf_num==0 && local_vf_num==1830 && local_vf_active==1) `fifo_error_check(1830)
              else if (local_pf_num==0 && local_vf_num==1831 && local_vf_active==1) `fifo_error_check(1831)
              else if (local_pf_num==0 && local_vf_num==1832 && local_vf_active==1) `fifo_error_check(1832)
              else if (local_pf_num==0 && local_vf_num==1833 && local_vf_active==1) `fifo_error_check(1833)
              else if (local_pf_num==0 && local_vf_num==1834 && local_vf_active==1) `fifo_error_check(1834)
              else if (local_pf_num==0 && local_vf_num==1835 && local_vf_active==1) `fifo_error_check(1835)
              else if (local_pf_num==0 && local_vf_num==1836 && local_vf_active==1) `fifo_error_check(1836)
              else if (local_pf_num==0 && local_vf_num==1837 && local_vf_active==1) `fifo_error_check(1837)
              else if (local_pf_num==0 && local_vf_num==1838 && local_vf_active==1) `fifo_error_check(1838)
              else if (local_pf_num==0 && local_vf_num==1839 && local_vf_active==1) `fifo_error_check(1839)
              else if (local_pf_num==0 && local_vf_num==1840 && local_vf_active==1) `fifo_error_check(1840)
              else if (local_pf_num==0 && local_vf_num==1841 && local_vf_active==1) `fifo_error_check(1841)
              else if (local_pf_num==0 && local_vf_num==1842 && local_vf_active==1) `fifo_error_check(1842)
              else if (local_pf_num==0 && local_vf_num==1843 && local_vf_active==1) `fifo_error_check(1843)
              else if (local_pf_num==0 && local_vf_num==1844 && local_vf_active==1) `fifo_error_check(1844)
              else if (local_pf_num==0 && local_vf_num==1845 && local_vf_active==1) `fifo_error_check(1845)
              else if (local_pf_num==0 && local_vf_num==1846 && local_vf_active==1) `fifo_error_check(1846)
              else if (local_pf_num==0 && local_vf_num==1847 && local_vf_active==1) `fifo_error_check(1847)
              else if (local_pf_num==0 && local_vf_num==1848 && local_vf_active==1) `fifo_error_check(1848)
              else if (local_pf_num==0 && local_vf_num==1849 && local_vf_active==1) `fifo_error_check(1849)
              else if (local_pf_num==0 && local_vf_num==1850 && local_vf_active==1) `fifo_error_check(1850)
              else if (local_pf_num==0 && local_vf_num==1851 && local_vf_active==1) `fifo_error_check(1851)
              else if (local_pf_num==0 && local_vf_num==1852 && local_vf_active==1) `fifo_error_check(1852)
              else if (local_pf_num==0 && local_vf_num==1853 && local_vf_active==1) `fifo_error_check(1853)
              else if (local_pf_num==0 && local_vf_num==1854 && local_vf_active==1) `fifo_error_check(1854)
              else if (local_pf_num==0 && local_vf_num==1855 && local_vf_active==1) `fifo_error_check(1855)
              else if (local_pf_num==0 && local_vf_num==1856 && local_vf_active==1) `fifo_error_check(1856)
              else if (local_pf_num==0 && local_vf_num==1857 && local_vf_active==1) `fifo_error_check(1857)
              else if (local_pf_num==0 && local_vf_num==1858 && local_vf_active==1) `fifo_error_check(1858)
              else if (local_pf_num==0 && local_vf_num==1859 && local_vf_active==1) `fifo_error_check(1859)
              else if (local_pf_num==0 && local_vf_num==1860 && local_vf_active==1) `fifo_error_check(1860)
              else if (local_pf_num==0 && local_vf_num==1861 && local_vf_active==1) `fifo_error_check(1861)
              else if (local_pf_num==0 && local_vf_num==1862 && local_vf_active==1) `fifo_error_check(1862)
              else if (local_pf_num==0 && local_vf_num==1863 && local_vf_active==1) `fifo_error_check(1863)
              else if (local_pf_num==0 && local_vf_num==1864 && local_vf_active==1) `fifo_error_check(1864)
              else if (local_pf_num==0 && local_vf_num==1865 && local_vf_active==1) `fifo_error_check(1865)
              else if (local_pf_num==0 && local_vf_num==1866 && local_vf_active==1) `fifo_error_check(1866)
              else if (local_pf_num==0 && local_vf_num==1867 && local_vf_active==1) `fifo_error_check(1867)
              else if (local_pf_num==0 && local_vf_num==1868 && local_vf_active==1) `fifo_error_check(1868)
              else if (local_pf_num==0 && local_vf_num==1869 && local_vf_active==1) `fifo_error_check(1869)
              else if (local_pf_num==0 && local_vf_num==1870 && local_vf_active==1) `fifo_error_check(1870)
              else if (local_pf_num==0 && local_vf_num==1871 && local_vf_active==1) `fifo_error_check(1871)
              else if (local_pf_num==0 && local_vf_num==1872 && local_vf_active==1) `fifo_error_check(1872)
              else if (local_pf_num==0 && local_vf_num==1873 && local_vf_active==1) `fifo_error_check(1873)
              else if (local_pf_num==0 && local_vf_num==1874 && local_vf_active==1) `fifo_error_check(1874)
              else if (local_pf_num==0 && local_vf_num==1875 && local_vf_active==1) `fifo_error_check(1875)
              else if (local_pf_num==0 && local_vf_num==1876 && local_vf_active==1) `fifo_error_check(1876)
              else if (local_pf_num==0 && local_vf_num==1877 && local_vf_active==1) `fifo_error_check(1877)
              else if (local_pf_num==0 && local_vf_num==1878 && local_vf_active==1) `fifo_error_check(1878)
              else if (local_pf_num==0 && local_vf_num==1879 && local_vf_active==1) `fifo_error_check(1879)
              else if (local_pf_num==0 && local_vf_num==1880 && local_vf_active==1) `fifo_error_check(1880)
              else if (local_pf_num==0 && local_vf_num==1881 && local_vf_active==1) `fifo_error_check(1881)
              else if (local_pf_num==0 && local_vf_num==1882 && local_vf_active==1) `fifo_error_check(1882)
              else if (local_pf_num==0 && local_vf_num==1883 && local_vf_active==1) `fifo_error_check(1883)
              else if (local_pf_num==0 && local_vf_num==1884 && local_vf_active==1) `fifo_error_check(1884)
              else if (local_pf_num==0 && local_vf_num==1885 && local_vf_active==1) `fifo_error_check(1885)
              else if (local_pf_num==0 && local_vf_num==1886 && local_vf_active==1) `fifo_error_check(1886)
              else if (local_pf_num==0 && local_vf_num==1887 && local_vf_active==1) `fifo_error_check(1887)
              else if (local_pf_num==0 && local_vf_num==1888 && local_vf_active==1) `fifo_error_check(1888)
              else if (local_pf_num==0 && local_vf_num==1889 && local_vf_active==1) `fifo_error_check(1889)
              else if (local_pf_num==0 && local_vf_num==1890 && local_vf_active==1) `fifo_error_check(1890)
              else if (local_pf_num==0 && local_vf_num==1891 && local_vf_active==1) `fifo_error_check(1891)
              else if (local_pf_num==0 && local_vf_num==1892 && local_vf_active==1) `fifo_error_check(1892)
              else if (local_pf_num==0 && local_vf_num==1893 && local_vf_active==1) `fifo_error_check(1893)
              else if (local_pf_num==0 && local_vf_num==1894 && local_vf_active==1) `fifo_error_check(1894)
              else if (local_pf_num==0 && local_vf_num==1895 && local_vf_active==1) `fifo_error_check(1895)
              else if (local_pf_num==0 && local_vf_num==1896 && local_vf_active==1) `fifo_error_check(1896)
              else if (local_pf_num==0 && local_vf_num==1897 && local_vf_active==1) `fifo_error_check(1897)
              else if (local_pf_num==0 && local_vf_num==1898 && local_vf_active==1) `fifo_error_check(1898)
              else if (local_pf_num==0 && local_vf_num==1899 && local_vf_active==1) `fifo_error_check(1899)
              else if (local_pf_num==0 && local_vf_num==1900 && local_vf_active==1) `fifo_error_check(1900)
              else if (local_pf_num==0 && local_vf_num==1901 && local_vf_active==1) `fifo_error_check(1901)
              else if (local_pf_num==0 && local_vf_num==1902 && local_vf_active==1) `fifo_error_check(1902)
              else if (local_pf_num==0 && local_vf_num==1903 && local_vf_active==1) `fifo_error_check(1903)
              else if (local_pf_num==0 && local_vf_num==1904 && local_vf_active==1) `fifo_error_check(1904)
              else if (local_pf_num==0 && local_vf_num==1905 && local_vf_active==1) `fifo_error_check(1905)
              else if (local_pf_num==0 && local_vf_num==1906 && local_vf_active==1) `fifo_error_check(1906)
              else if (local_pf_num==0 && local_vf_num==1907 && local_vf_active==1) `fifo_error_check(1907)
              else if (local_pf_num==0 && local_vf_num==1908 && local_vf_active==1) `fifo_error_check(1908)
              else if (local_pf_num==0 && local_vf_num==1909 && local_vf_active==1) `fifo_error_check(1909)
              else if (local_pf_num==0 && local_vf_num==1910 && local_vf_active==1) `fifo_error_check(1910)
              else if (local_pf_num==0 && local_vf_num==1911 && local_vf_active==1) `fifo_error_check(1911)
              else if (local_pf_num==0 && local_vf_num==1912 && local_vf_active==1) `fifo_error_check(1912)
              else if (local_pf_num==0 && local_vf_num==1913 && local_vf_active==1) `fifo_error_check(1913)
              else if (local_pf_num==0 && local_vf_num==1914 && local_vf_active==1) `fifo_error_check(1914)
              else if (local_pf_num==0 && local_vf_num==1915 && local_vf_active==1) `fifo_error_check(1915)
              else if (local_pf_num==0 && local_vf_num==1916 && local_vf_active==1) `fifo_error_check(1916)
              else if (local_pf_num==0 && local_vf_num==1917 && local_vf_active==1) `fifo_error_check(1917)
              else if (local_pf_num==0 && local_vf_num==1918 && local_vf_active==1) `fifo_error_check(1918)
              else if (local_pf_num==0 && local_vf_num==1919 && local_vf_active==1) `fifo_error_check(1919)
              else if (local_pf_num==0 && local_vf_num==1920 && local_vf_active==1) `fifo_error_check(1920)
              else if (local_pf_num==0 && local_vf_num==1921 && local_vf_active==1) `fifo_error_check(1921)
              else if (local_pf_num==0 && local_vf_num==1922 && local_vf_active==1) `fifo_error_check(1922)
              else if (local_pf_num==0 && local_vf_num==1923 && local_vf_active==1) `fifo_error_check(1923)
              else if (local_pf_num==0 && local_vf_num==1924 && local_vf_active==1) `fifo_error_check(1924)
              else if (local_pf_num==0 && local_vf_num==1925 && local_vf_active==1) `fifo_error_check(1925)
              else if (local_pf_num==0 && local_vf_num==1926 && local_vf_active==1) `fifo_error_check(1926)
              else if (local_pf_num==0 && local_vf_num==1927 && local_vf_active==1) `fifo_error_check(1927)
              else if (local_pf_num==0 && local_vf_num==1928 && local_vf_active==1) `fifo_error_check(1928)
              else if (local_pf_num==0 && local_vf_num==1929 && local_vf_active==1) `fifo_error_check(1929)
              else if (local_pf_num==0 && local_vf_num==1930 && local_vf_active==1) `fifo_error_check(1930)
              else if (local_pf_num==0 && local_vf_num==1931 && local_vf_active==1) `fifo_error_check(1931)
              else if (local_pf_num==0 && local_vf_num==1932 && local_vf_active==1) `fifo_error_check(1932)
              else if (local_pf_num==0 && local_vf_num==1933 && local_vf_active==1) `fifo_error_check(1933)
              else if (local_pf_num==0 && local_vf_num==1934 && local_vf_active==1) `fifo_error_check(1934)
              else if (local_pf_num==0 && local_vf_num==1935 && local_vf_active==1) `fifo_error_check(1935)
              else if (local_pf_num==0 && local_vf_num==1936 && local_vf_active==1) `fifo_error_check(1936)
              else if (local_pf_num==0 && local_vf_num==1937 && local_vf_active==1) `fifo_error_check(1937)
              else if (local_pf_num==0 && local_vf_num==1938 && local_vf_active==1) `fifo_error_check(1938)
              else if (local_pf_num==0 && local_vf_num==1939 && local_vf_active==1) `fifo_error_check(1939)
              else if (local_pf_num==0 && local_vf_num==1940 && local_vf_active==1) `fifo_error_check(1940)
              else if (local_pf_num==0 && local_vf_num==1941 && local_vf_active==1) `fifo_error_check(1941)
              else if (local_pf_num==0 && local_vf_num==1942 && local_vf_active==1) `fifo_error_check(1942)
              else if (local_pf_num==0 && local_vf_num==1943 && local_vf_active==1) `fifo_error_check(1943)
              else if (local_pf_num==0 && local_vf_num==1944 && local_vf_active==1) `fifo_error_check(1944)
              else if (local_pf_num==0 && local_vf_num==1945 && local_vf_active==1) `fifo_error_check(1945)
              else if (local_pf_num==0 && local_vf_num==1946 && local_vf_active==1) `fifo_error_check(1946)
              else if (local_pf_num==0 && local_vf_num==1947 && local_vf_active==1) `fifo_error_check(1947)
              else if (local_pf_num==0 && local_vf_num==1948 && local_vf_active==1) `fifo_error_check(1948)
              else if (local_pf_num==0 && local_vf_num==1949 && local_vf_active==1) `fifo_error_check(1949)
              else if (local_pf_num==0 && local_vf_num==1950 && local_vf_active==1) `fifo_error_check(1950)
              else if (local_pf_num==0 && local_vf_num==1951 && local_vf_active==1) `fifo_error_check(1951)
              else if (local_pf_num==0 && local_vf_num==1952 && local_vf_active==1) `fifo_error_check(1952)
              else if (local_pf_num==0 && local_vf_num==1953 && local_vf_active==1) `fifo_error_check(1953)
              else if (local_pf_num==0 && local_vf_num==1954 && local_vf_active==1) `fifo_error_check(1954)
              else if (local_pf_num==0 && local_vf_num==1955 && local_vf_active==1) `fifo_error_check(1955)
              else if (local_pf_num==0 && local_vf_num==1956 && local_vf_active==1) `fifo_error_check(1956)
              else if (local_pf_num==0 && local_vf_num==1957 && local_vf_active==1) `fifo_error_check(1957)
              else if (local_pf_num==0 && local_vf_num==1958 && local_vf_active==1) `fifo_error_check(1958)
              else if (local_pf_num==0 && local_vf_num==1959 && local_vf_active==1) `fifo_error_check(1959)
              else if (local_pf_num==0 && local_vf_num==1960 && local_vf_active==1) `fifo_error_check(1960)
              else if (local_pf_num==0 && local_vf_num==1961 && local_vf_active==1) `fifo_error_check(1961)
              else if (local_pf_num==0 && local_vf_num==1962 && local_vf_active==1) `fifo_error_check(1962)
              else if (local_pf_num==0 && local_vf_num==1963 && local_vf_active==1) `fifo_error_check(1963)
              else if (local_pf_num==0 && local_vf_num==1964 && local_vf_active==1) `fifo_error_check(1964)
              else if (local_pf_num==0 && local_vf_num==1965 && local_vf_active==1) `fifo_error_check(1965)
              else if (local_pf_num==0 && local_vf_num==1966 && local_vf_active==1) `fifo_error_check(1966)
              else if (local_pf_num==0 && local_vf_num==1967 && local_vf_active==1) `fifo_error_check(1967)
              else if (local_pf_num==0 && local_vf_num==1968 && local_vf_active==1) `fifo_error_check(1968)
              else if (local_pf_num==0 && local_vf_num==1969 && local_vf_active==1) `fifo_error_check(1969)
              else if (local_pf_num==0 && local_vf_num==1970 && local_vf_active==1) `fifo_error_check(1970)
              else if (local_pf_num==0 && local_vf_num==1971 && local_vf_active==1) `fifo_error_check(1971)
              else if (local_pf_num==0 && local_vf_num==1972 && local_vf_active==1) `fifo_error_check(1972)
              else if (local_pf_num==0 && local_vf_num==1973 && local_vf_active==1) `fifo_error_check(1973)
              else if (local_pf_num==0 && local_vf_num==1974 && local_vf_active==1) `fifo_error_check(1974)
              else if (local_pf_num==0 && local_vf_num==1975 && local_vf_active==1) `fifo_error_check(1975)
              else if (local_pf_num==0 && local_vf_num==1976 && local_vf_active==1) `fifo_error_check(1976)
              else if (local_pf_num==0 && local_vf_num==1977 && local_vf_active==1) `fifo_error_check(1977)
              else if (local_pf_num==0 && local_vf_num==1978 && local_vf_active==1) `fifo_error_check(1978)
              else if (local_pf_num==0 && local_vf_num==1979 && local_vf_active==1) `fifo_error_check(1979)
              else if (local_pf_num==0 && local_vf_num==1980 && local_vf_active==1) `fifo_error_check(1980)
              else if (local_pf_num==0 && local_vf_num==1981 && local_vf_active==1) `fifo_error_check(1981)
              else if (local_pf_num==0 && local_vf_num==1982 && local_vf_active==1) `fifo_error_check(1982)
              else if (local_pf_num==0 && local_vf_num==1983 && local_vf_active==1) `fifo_error_check(1983)
              else if (local_pf_num==0 && local_vf_num==1984 && local_vf_active==1) `fifo_error_check(1984)
              else if (local_pf_num==0 && local_vf_num==1985 && local_vf_active==1) `fifo_error_check(1985)
              else if (local_pf_num==0 && local_vf_num==1986 && local_vf_active==1) `fifo_error_check(1986)
              else if (local_pf_num==0 && local_vf_num==1987 && local_vf_active==1) `fifo_error_check(1987)
              else if (local_pf_num==0 && local_vf_num==1988 && local_vf_active==1) `fifo_error_check(1988)
              else if (local_pf_num==0 && local_vf_num==1989 && local_vf_active==1) `fifo_error_check(1989)
              else if (local_pf_num==0 && local_vf_num==1990 && local_vf_active==1) `fifo_error_check(1990)
              else if (local_pf_num==0 && local_vf_num==1991 && local_vf_active==1) `fifo_error_check(1991)
              else if (local_pf_num==0 && local_vf_num==1992 && local_vf_active==1) `fifo_error_check(1992)
              else if (local_pf_num==0 && local_vf_num==1993 && local_vf_active==1) `fifo_error_check(1993)
              else if (local_pf_num==0 && local_vf_num==1994 && local_vf_active==1) `fifo_error_check(1994)
              else if (local_pf_num==0 && local_vf_num==1995 && local_vf_active==1) `fifo_error_check(1995)
              else if (local_pf_num==0 && local_vf_num==1996 && local_vf_active==1) `fifo_error_check(1996)
              else if (local_pf_num==0 && local_vf_num==1997 && local_vf_active==1) `fifo_error_check(1997)
              else if (local_pf_num==0 && local_vf_num==1998 && local_vf_active==1) `fifo_error_check(1998)
              else if (local_pf_num==0 && local_vf_num==1999 && local_vf_active==1) `fifo_error_check(1999)
              else if (local_pf_num==0 && local_vf_num==2000 && local_vf_active==1) `fifo_error_check(2000)
              else if (local_pf_num==0 && local_vf_num==2001 && local_vf_active==1) `fifo_error_check(2001)
              else if (local_pf_num==0 && local_vf_num==2002 && local_vf_active==1) `fifo_error_check(2002)
              else if (local_pf_num==0 && local_vf_num==2003 && local_vf_active==1) `fifo_error_check(2003)
              else if (local_pf_num==0 && local_vf_num==2004 && local_vf_active==1) `fifo_error_check(2004)
              else if (local_pf_num==0 && local_vf_num==2005 && local_vf_active==1) `fifo_error_check(2005)
              else if (local_pf_num==0 && local_vf_num==2006 && local_vf_active==1) `fifo_error_check(2006)
              else if (local_pf_num==0 && local_vf_num==2007 && local_vf_active==1) `fifo_error_check(2007)
              else if (local_pf_num==0 && local_vf_num==2008 && local_vf_active==1) `fifo_error_check(2008)
              else if (local_pf_num==0 && local_vf_num==2009 && local_vf_active==1) `fifo_error_check(2009)
              else if (local_pf_num==0 && local_vf_num==2010 && local_vf_active==1) `fifo_error_check(2010)
              else if (local_pf_num==0 && local_vf_num==2011 && local_vf_active==1) `fifo_error_check(2011)
              else if (local_pf_num==0 && local_vf_num==2012 && local_vf_active==1) `fifo_error_check(2012)
              else if (local_pf_num==0 && local_vf_num==2013 && local_vf_active==1) `fifo_error_check(2013)
              else if (local_pf_num==0 && local_vf_num==2014 && local_vf_active==1) `fifo_error_check(2014)
              else if (local_pf_num==0 && local_vf_num==2015 && local_vf_active==1) `fifo_error_check(2015)
              else if (local_pf_num==0 && local_vf_num==2016 && local_vf_active==1) `fifo_error_check(2016)
              else if (local_pf_num==0 && local_vf_num==2017 && local_vf_active==1) `fifo_error_check(2017)
              else if (local_pf_num==0 && local_vf_num==2018 && local_vf_active==1) `fifo_error_check(2018)
              else if (local_pf_num==0 && local_vf_num==2019 && local_vf_active==1) `fifo_error_check(2019)
              else if (local_pf_num==0 && local_vf_num==2020 && local_vf_active==1) `fifo_error_check(2020)
              else if (local_pf_num==0 && local_vf_num==2021 && local_vf_active==1) `fifo_error_check(2021)
              else if (local_pf_num==0 && local_vf_num==2022 && local_vf_active==1) `fifo_error_check(2022)
              else if (local_pf_num==0 && local_vf_num==2023 && local_vf_active==1) `fifo_error_check(2023)
              else if (local_pf_num==0 && local_vf_num==2024 && local_vf_active==1) `fifo_error_check(2024)
              else if (local_pf_num==0 && local_vf_num==2025 && local_vf_active==1) `fifo_error_check(2025)
              else if (local_pf_num==0 && local_vf_num==2026 && local_vf_active==1) `fifo_error_check(2026)
              else if (local_pf_num==0 && local_vf_num==2027 && local_vf_active==1) `fifo_error_check(2027)
              else if (local_pf_num==0 && local_vf_num==2028 && local_vf_active==1) `fifo_error_check(2028)
              else if (local_pf_num==0 && local_vf_num==2029 && local_vf_active==1) `fifo_error_check(2029)
              else if (local_pf_num==0 && local_vf_num==2030 && local_vf_active==1) `fifo_error_check(2030)
              else if (local_pf_num==0 && local_vf_num==2031 && local_vf_active==1) `fifo_error_check(2031)
              else if (local_pf_num==0 && local_vf_num==2032 && local_vf_active==1) `fifo_error_check(2032)
              else if (local_pf_num==0 && local_vf_num==2033 && local_vf_active==1) `fifo_error_check(2033)
              else if (local_pf_num==0 && local_vf_num==2034 && local_vf_active==1) `fifo_error_check(2034)
              else if (local_pf_num==0 && local_vf_num==2035 && local_vf_active==1) `fifo_error_check(2035)
              else if (local_pf_num==0 && local_vf_num==2036 && local_vf_active==1) `fifo_error_check(2036)
              else if (local_pf_num==0 && local_vf_num==2037 && local_vf_active==1) `fifo_error_check(2037)
              else if (local_pf_num==0 && local_vf_num==2038 && local_vf_active==1) `fifo_error_check(2038)
              else if (local_pf_num==0 && local_vf_num==2039 && local_vf_active==1) `fifo_error_check(2039)
              else if (local_pf_num==0 && local_vf_num==2040 && local_vf_active==1) `fifo_error_check(2040)
              else if (local_pf_num==0 && local_vf_num==2041 && local_vf_active==1) `fifo_error_check(2041)
              else if (local_pf_num==0 && local_vf_num==2042 && local_vf_active==1) `fifo_error_check(2042)
              else if (local_pf_num==0 && local_vf_num==2043 && local_vf_active==1) `fifo_error_check(2043)
              else if (local_pf_num==0 && local_vf_num==2044 && local_vf_active==1) `fifo_error_check(2044)
              else if (local_pf_num==0 && local_vf_num==2045 && local_vf_active==1) `fifo_error_check(2045)
              else if (local_pf_num==0 && local_vf_num==2046 && local_vf_active==1) `fifo_error_check(2046)
              else if (local_pf_num==0 && local_vf_num==2047 && local_vf_active==1) `fifo_error_check(2047)
              `endif 

        fork
          begin
              `ifdef TB_CONFIG_1
              if (local_pf_num==0 && local_vf_num ==0 && local_vf_active==0) 
                 `toggle_tready(0)   
              else if (local_pf_num==1 && local_vf_num==0 && local_vf_active==0) 
                `toggle_tready(1)                     
              else if (local_pf_num==2 && local_vf_num==0 && local_vf_active==0) 
                 `toggle_tready(2)                    
              else if (local_pf_num==3 && local_vf_num==0 && local_vf_active==0) 
                  `toggle_tready(3)                   
              else if (local_pf_num==4 && local_vf_num==0 && local_vf_active==0) 
                  `toggle_tready(4)                                  
              else if (local_pf_num==5 && local_vf_num==0 && local_vf_active==0) 
                   `toggle_tready(5)                                 
              else if (local_pf_num==6 && local_vf_num==0 && local_vf_active==0) 
                   `toggle_tready(6)                  
              else if (local_pf_num==7 && local_vf_num==0 && local_vf_active==0) 
                    `toggle_tready(7)                    
              else if (local_pf_num==0 && local_vf_num==0 && local_vf_active==1) 
                    `toggle_tready(8)                    
              else if (local_pf_num==1 && local_vf_num==0 && local_vf_active==1) 
                    `toggle_tready(9)     
              else if (local_pf_num==2 && local_vf_num==0 && local_vf_active==1) 
                   `toggle_tready(10)                    
              else if (local_pf_num==3 && local_vf_num==0 && local_vf_active==1) 
                   `toggle_tready(11)                    
              else if (local_pf_num==4 && local_vf_num==0 && local_vf_active==1) 
                   `toggle_tready(12)     
              else if (local_pf_num==5 && local_vf_num==0 && local_vf_active==1) 
                   `toggle_tready(13)                    
              else if (local_pf_num==6 && local_vf_num==0 && local_vf_active==1) 
                   `toggle_tready(14)                    
              else if (local_pf_num==7 && local_vf_num==0 && local_vf_active==1) 
                    `toggle_tready(15)

              `elsif TB_CONFIG_2
              if (local_pf_num==0 && local_vf_num ==0 && local_vf_active==0) 
                 `toggle_tready(0)   
              else if (local_pf_num==1 && local_vf_num==0 && local_vf_active==0) 
                `toggle_tready(1)                     
              else if (local_pf_num==2 && local_vf_num==0 && local_vf_active==0) 
                 `toggle_tready(2)                    
              else if (local_pf_num==3 && local_vf_num==0 && local_vf_active==0) 
                  `toggle_tready(3)                   
              else if (local_pf_num==4 && local_vf_num==0 && local_vf_active==0) 
                  `toggle_tready(4)                                  
              else if (local_pf_num==5 && local_vf_num==0 && local_vf_active==0) 
                   `toggle_tready(5)                                 
              else if (local_pf_num==6 && local_vf_num==0 && local_vf_active==0) 
                   `toggle_tready(6)                  
              else if (local_pf_num==7 && local_vf_num==0 && local_vf_active==0) 
                    `toggle_tready(7)                    
              else if (local_pf_num==0 && local_vf_num==0 && local_vf_active==1) 
                    `toggle_tready(8)                    
              else if (local_pf_num==1 && local_vf_num==0 && local_vf_active==1) 
                    `toggle_tready(9)     
              else if (local_pf_num==2 && local_vf_num==0 && local_vf_active==1) 
                   `toggle_tready(10)                    
              else if (local_pf_num==3 && local_vf_num==0 && local_vf_active==1) 
                   `toggle_tready(11)                    
              else if (local_pf_num==4 && local_vf_num==0 && local_vf_active==1) 
                   `toggle_tready(12)     
              else if (local_pf_num==5 && local_vf_num==0 && local_vf_active==1) 
                   `toggle_tready(13)                    
              else if (local_pf_num==6 && local_vf_num==0 && local_vf_active==1) 
                   `toggle_tready(14)                    
              else if (local_pf_num==7 && local_vf_num==0 && local_vf_active==1) 
                    `toggle_tready(15)
              else if (local_pf_num==0 && local_vf_num=='h7ff && local_vf_active==1) 
                    `toggle_tready(16)                                             
              else if (local_pf_num==1 && local_vf_num=='h7ff && local_vf_active==1) 
                    `toggle_tready(17)                                             
              else if (local_pf_num==2 && local_vf_num=='h7ff && local_vf_active==1) 
                   `toggle_tready(18)                                              
              else if (local_pf_num==3 && local_vf_num=='h7ff && local_vf_active==1) 
                   `toggle_tready(19)                                              
              else if (local_pf_num==4 && local_vf_num=='h7ff && local_vf_active==1) 
                   `toggle_tready(20)                                             
              else if (local_pf_num==5 && local_vf_num=='h7ff && local_vf_active==1) 
                   `toggle_tready(21)                                          
              else if (local_pf_num==6 && local_vf_num=='h7ff && local_vf_active==1) 
                   `toggle_tready(22)
              else if (local_pf_num==7 && local_vf_num=='h7ff && local_vf_active==1) 
                    `toggle_tready(23)

              `elsif TB_CONFIG_3
              if (local_pf_num==0 && local_vf_num ==0 && local_vf_active==0) 
                 `toggle_tready(0)   
              else if (local_pf_num==1 && local_vf_num==0 && local_vf_active==0) 
                `toggle_tready(1)                     
              else if (local_pf_num==2 && local_vf_num==0 && local_vf_active==0) 
                 `toggle_tready(2)                    
              else if (local_pf_num==3 && local_vf_num==0 && local_vf_active==0) 
                  `toggle_tready(3)                   
              else if (local_pf_num==4 && local_vf_num==0 && local_vf_active==0) 
                  `toggle_tready(4)                                  
              else if (local_pf_num==5 && local_vf_num==0 && local_vf_active==0) 
                   `toggle_tready(5)                                 
              else if (local_pf_num==6 && local_vf_num==0 && local_vf_active==0) 
                   `toggle_tready(6)                  
              else if (local_pf_num==7 && local_vf_num==0 && local_vf_active==0) 
                    `toggle_tready(7)                    
              else if (local_pf_num==0 && local_vf_num==0 && local_vf_active==1) 
                    `toggle_tready(8)                    
              else if (local_pf_num==1 && local_vf_num==0 && local_vf_active==1) 
                    `toggle_tready(9)     
              else if (local_pf_num==2 && local_vf_num==0 && local_vf_active==1) 
                   `toggle_tready(10)                    
              else if (local_pf_num==3 && local_vf_num==0 && local_vf_active==1) 
                   `toggle_tready(11)                    
              else if (local_pf_num==4 && local_vf_num==0 && local_vf_active==1) 
                   `toggle_tready(12)     
              else if (local_pf_num==5 && local_vf_num==0 && local_vf_active==1) 
                   `toggle_tready(13)                    
              else if (local_pf_num==6 && local_vf_num==0 && local_vf_active==1) 
                   `toggle_tready(14)                    
              else if (local_pf_num==7 && local_vf_num==0 && local_vf_active==1) 
                    `toggle_tready(15)
              else if (local_pf_num==0 && local_vf_num=='h7ff && local_vf_active==1) 
                    `toggle_tready(16)                                             
              else if (local_pf_num==1 && local_vf_num=='h7ff && local_vf_active==1) 
                    `toggle_tready(17)                                             
              else if (local_pf_num==2 && local_vf_num=='h7ff && local_vf_active==1) 
                   `toggle_tready(18)                                              
              else if (local_pf_num==3 && local_vf_num=='h7ff && local_vf_active==1) 
                   `toggle_tready(19)                                              
              else if (local_pf_num==4 && local_vf_num=='h7ff && local_vf_active==1) 
                   `toggle_tready(20)                                             
              else if (local_pf_num==5 && local_vf_num=='h7ff && local_vf_active==1) 
                   `toggle_tready(21)                                          
              else if (local_pf_num==6 && local_vf_num=='h7ff && local_vf_active==1) 
                   `toggle_tready(22)
              else if (local_pf_num==7 && local_vf_num=='h7ff && local_vf_active==1) 
                    `toggle_tready(23)
              else if (local_pf_num==0 && local_vf_num==`RANDOM_VF && local_vf_active==1) 
                    `toggle_tready(24)                                        
              else if (local_pf_num==1 && local_vf_num==`RANDOM_VF && local_vf_active==1) 
                    `toggle_tready(25)                                        
              else if (local_pf_num==2 && local_vf_num==`RANDOM_VF && local_vf_active==1) 
                   `toggle_tready(26)                                         
              else if (local_pf_num==3 && local_vf_num==`RANDOM_VF && local_vf_active==1) 
                   `toggle_tready(27)                                         
              else if (local_pf_num==4 && local_vf_num==`RANDOM_VF && local_vf_active==1) 
                   `toggle_tready(28)                                        
              else if (local_pf_num==5 && local_vf_num==`RANDOM_VF && local_vf_active==1) 
                   `toggle_tready(29)                                     
              else if (local_pf_num==6 && local_vf_num==`RANDOM_VF && local_vf_active==1) 
                   `toggle_tready(30)
              else if (local_pf_num==7 && local_vf_num==`RANDOM_VF && local_vf_active==1) 
                    `toggle_tready(31)
              `elsif TB_CONFIG_4
              if (local_pf_num==0 && local_vf_num ==0 && local_vf_active==1) `toggle_tready(0)   
              else if (local_pf_num==0 && local_vf_num ==1 && local_vf_active==1) `toggle_tready(1)   
              else if (local_pf_num==0 && local_vf_num ==2 && local_vf_active==1) `toggle_tready(2)   
              else if (local_pf_num==0 && local_vf_num ==3 && local_vf_active==1) `toggle_tready(3)   
              else if (local_pf_num==0 && local_vf_num ==4 && local_vf_active==1) `toggle_tready(4)   
              else if (local_pf_num==0 && local_vf_num ==5 && local_vf_active==1) `toggle_tready(5)   
              else if (local_pf_num==0 && local_vf_num ==6 && local_vf_active==1) `toggle_tready(6)   
              else if (local_pf_num==0 && local_vf_num ==7 && local_vf_active==1) `toggle_tready(7)   
              else if (local_pf_num==0 && local_vf_num ==8 && local_vf_active==1) `toggle_tready(8)   
              else if (local_pf_num==0 && local_vf_num ==9 && local_vf_active==1) `toggle_tready(9)   
              else if (local_pf_num==0 && local_vf_num ==10 && local_vf_active==1) `toggle_tready(10)   
              else if (local_pf_num==0 && local_vf_num ==11 && local_vf_active==1) `toggle_tready(11)   
              else if (local_pf_num==0 && local_vf_num ==12 && local_vf_active==1) `toggle_tready(12)   
              else if (local_pf_num==0 && local_vf_num ==13 && local_vf_active==1) `toggle_tready(13)   
              else if (local_pf_num==0 && local_vf_num ==14 && local_vf_active==1) `toggle_tready(14)   
              else if (local_pf_num==0 && local_vf_num ==15 && local_vf_active==1) `toggle_tready(15)   
              else if (local_pf_num==0 && local_vf_num ==16 && local_vf_active==1) `toggle_tready(16)   
              else if (local_pf_num==0 && local_vf_num ==17 && local_vf_active==1) `toggle_tready(17)   
              else if (local_pf_num==0 && local_vf_num ==18 && local_vf_active==1) `toggle_tready(18)   
              else if (local_pf_num==0 && local_vf_num ==19 && local_vf_active==1) `toggle_tready(19)   
              else if (local_pf_num==0 && local_vf_num ==20 && local_vf_active==1) `toggle_tready(20)   
              else if (local_pf_num==0 && local_vf_num ==21 && local_vf_active==1) `toggle_tready(21)   
              else if (local_pf_num==0 && local_vf_num ==22 && local_vf_active==1) `toggle_tready(22)   
              else if (local_pf_num==0 && local_vf_num ==23 && local_vf_active==1) `toggle_tready(23)   
              else if (local_pf_num==0 && local_vf_num ==24 && local_vf_active==1) `toggle_tready(24)   
              else if (local_pf_num==0 && local_vf_num ==25 && local_vf_active==1) `toggle_tready(25)   
              else if (local_pf_num==0 && local_vf_num ==26 && local_vf_active==1) `toggle_tready(26)   
              else if (local_pf_num==0 && local_vf_num ==27 && local_vf_active==1) `toggle_tready(27)   
              else if (local_pf_num==0 && local_vf_num ==28 && local_vf_active==1) `toggle_tready(28)   
              else if (local_pf_num==0 && local_vf_num ==29 && local_vf_active==1) `toggle_tready(29)   
              else if (local_pf_num==0 && local_vf_num ==30 && local_vf_active==1) `toggle_tready(30)   
              else if (local_pf_num==0 && local_vf_num ==31 && local_vf_active==1) `toggle_tready(31)   
              else if (local_pf_num==0 && local_vf_num ==32 && local_vf_active==1) `toggle_tready(32)   
              else if (local_pf_num==0 && local_vf_num ==33 && local_vf_active==1) `toggle_tready(33)   
              else if (local_pf_num==0 && local_vf_num ==34 && local_vf_active==1) `toggle_tready(34)   
              else if (local_pf_num==0 && local_vf_num ==35 && local_vf_active==1) `toggle_tready(35)   
              else if (local_pf_num==0 && local_vf_num ==36 && local_vf_active==1) `toggle_tready(36)   
              else if (local_pf_num==0 && local_vf_num ==37 && local_vf_active==1) `toggle_tready(37)   
              else if (local_pf_num==0 && local_vf_num ==38 && local_vf_active==1) `toggle_tready(38)   
              else if (local_pf_num==0 && local_vf_num ==39 && local_vf_active==1) `toggle_tready(39)   
              else if (local_pf_num==0 && local_vf_num ==40 && local_vf_active==1) `toggle_tready(40)   
              else if (local_pf_num==0 && local_vf_num ==41 && local_vf_active==1) `toggle_tready(41)   
              else if (local_pf_num==0 && local_vf_num ==42 && local_vf_active==1) `toggle_tready(42)   
              else if (local_pf_num==0 && local_vf_num ==43 && local_vf_active==1) `toggle_tready(43)   
              else if (local_pf_num==0 && local_vf_num ==44 && local_vf_active==1) `toggle_tready(44)   
              else if (local_pf_num==0 && local_vf_num ==45 && local_vf_active==1) `toggle_tready(45)   
              else if (local_pf_num==0 && local_vf_num ==46 && local_vf_active==1) `toggle_tready(46)   
              else if (local_pf_num==0 && local_vf_num ==47 && local_vf_active==1) `toggle_tready(47)   
              else if (local_pf_num==0 && local_vf_num ==48 && local_vf_active==1) `toggle_tready(48)   
              else if (local_pf_num==0 && local_vf_num ==49 && local_vf_active==1) `toggle_tready(49)   
              else if (local_pf_num==0 && local_vf_num ==50 && local_vf_active==1) `toggle_tready(50)   
              else if (local_pf_num==0 && local_vf_num ==51 && local_vf_active==1) `toggle_tready(51)   
              else if (local_pf_num==0 && local_vf_num ==52 && local_vf_active==1) `toggle_tready(52)   
              else if (local_pf_num==0 && local_vf_num ==53 && local_vf_active==1) `toggle_tready(53)   
              else if (local_pf_num==0 && local_vf_num ==54 && local_vf_active==1) `toggle_tready(54)   
              else if (local_pf_num==0 && local_vf_num ==55 && local_vf_active==1) `toggle_tready(55)   
              else if (local_pf_num==0 && local_vf_num ==56 && local_vf_active==1) `toggle_tready(56)   
              else if (local_pf_num==0 && local_vf_num ==57 && local_vf_active==1) `toggle_tready(57)   
              else if (local_pf_num==0 && local_vf_num ==58 && local_vf_active==1) `toggle_tready(58)   
              else if (local_pf_num==0 && local_vf_num ==59 && local_vf_active==1) `toggle_tready(59)   
              else if (local_pf_num==0 && local_vf_num ==60 && local_vf_active==1) `toggle_tready(60)   
              else if (local_pf_num==0 && local_vf_num ==61 && local_vf_active==1) `toggle_tready(61)   
              else if (local_pf_num==0 && local_vf_num ==62 && local_vf_active==1) `toggle_tready(62)   
              else if (local_pf_num==0 && local_vf_num ==63 && local_vf_active==1) `toggle_tready(63)   
              else if (local_pf_num==0 && local_vf_num ==64 && local_vf_active==1) `toggle_tready(64)   
              else if (local_pf_num==0 && local_vf_num ==65 && local_vf_active==1) `toggle_tready(65)   
              else if (local_pf_num==0 && local_vf_num ==66 && local_vf_active==1) `toggle_tready(66)   
              else if (local_pf_num==0 && local_vf_num ==67 && local_vf_active==1) `toggle_tready(67)   
              else if (local_pf_num==0 && local_vf_num ==68 && local_vf_active==1) `toggle_tready(68)   
              else if (local_pf_num==0 && local_vf_num ==69 && local_vf_active==1) `toggle_tready(69)   
              else if (local_pf_num==0 && local_vf_num ==70 && local_vf_active==1) `toggle_tready(70)   
              else if (local_pf_num==0 && local_vf_num ==71 && local_vf_active==1) `toggle_tready(71)   
              else if (local_pf_num==0 && local_vf_num ==72 && local_vf_active==1) `toggle_tready(72)   
              else if (local_pf_num==0 && local_vf_num ==73 && local_vf_active==1) `toggle_tready(73)   
              else if (local_pf_num==0 && local_vf_num ==74 && local_vf_active==1) `toggle_tready(74)   
              else if (local_pf_num==0 && local_vf_num ==75 && local_vf_active==1) `toggle_tready(75)   
              else if (local_pf_num==0 && local_vf_num ==76 && local_vf_active==1) `toggle_tready(76)   
              else if (local_pf_num==0 && local_vf_num ==77 && local_vf_active==1) `toggle_tready(77)   
              else if (local_pf_num==0 && local_vf_num ==78 && local_vf_active==1) `toggle_tready(78)   
              else if (local_pf_num==0 && local_vf_num ==79 && local_vf_active==1) `toggle_tready(79)   
              else if (local_pf_num==0 && local_vf_num ==80 && local_vf_active==1) `toggle_tready(80)   
              else if (local_pf_num==0 && local_vf_num ==81 && local_vf_active==1) `toggle_tready(81)   
              else if (local_pf_num==0 && local_vf_num ==82 && local_vf_active==1) `toggle_tready(82)   
              else if (local_pf_num==0 && local_vf_num ==83 && local_vf_active==1) `toggle_tready(83)   
              else if (local_pf_num==0 && local_vf_num ==84 && local_vf_active==1) `toggle_tready(84)   
              else if (local_pf_num==0 && local_vf_num ==85 && local_vf_active==1) `toggle_tready(85)   
              else if (local_pf_num==0 && local_vf_num ==86 && local_vf_active==1) `toggle_tready(86)   
              else if (local_pf_num==0 && local_vf_num ==87 && local_vf_active==1) `toggle_tready(87)   
              else if (local_pf_num==0 && local_vf_num ==88 && local_vf_active==1) `toggle_tready(88)   
              else if (local_pf_num==0 && local_vf_num ==89 && local_vf_active==1) `toggle_tready(89)   
              else if (local_pf_num==0 && local_vf_num ==90 && local_vf_active==1) `toggle_tready(90)   
              else if (local_pf_num==0 && local_vf_num ==91 && local_vf_active==1) `toggle_tready(91)   
              else if (local_pf_num==0 && local_vf_num ==92 && local_vf_active==1) `toggle_tready(92)   
              else if (local_pf_num==0 && local_vf_num ==93 && local_vf_active==1) `toggle_tready(93)   
              else if (local_pf_num==0 && local_vf_num ==94 && local_vf_active==1) `toggle_tready(94)   
              else if (local_pf_num==0 && local_vf_num ==95 && local_vf_active==1) `toggle_tready(95)   
              else if (local_pf_num==0 && local_vf_num ==96 && local_vf_active==1) `toggle_tready(96)   
              else if (local_pf_num==0 && local_vf_num ==97 && local_vf_active==1) `toggle_tready(97)   
              else if (local_pf_num==0 && local_vf_num ==98 && local_vf_active==1) `toggle_tready(98)   
              else if (local_pf_num==0 && local_vf_num ==99 && local_vf_active==1) `toggle_tready(99)   
              else if (local_pf_num==0 && local_vf_num ==100 && local_vf_active==1) `toggle_tready(100)   
              else if (local_pf_num==0 && local_vf_num ==101 && local_vf_active==1) `toggle_tready(101)   
              else if (local_pf_num==0 && local_vf_num ==102 && local_vf_active==1) `toggle_tready(102)   
              else if (local_pf_num==0 && local_vf_num ==103 && local_vf_active==1) `toggle_tready(103)   
              else if (local_pf_num==0 && local_vf_num ==104 && local_vf_active==1) `toggle_tready(104)   
              else if (local_pf_num==0 && local_vf_num ==105 && local_vf_active==1) `toggle_tready(105)   
              else if (local_pf_num==0 && local_vf_num ==106 && local_vf_active==1) `toggle_tready(106)   
              else if (local_pf_num==0 && local_vf_num ==107 && local_vf_active==1) `toggle_tready(107)   
              else if (local_pf_num==0 && local_vf_num ==108 && local_vf_active==1) `toggle_tready(108)   
              else if (local_pf_num==0 && local_vf_num ==109 && local_vf_active==1) `toggle_tready(109)   
              else if (local_pf_num==0 && local_vf_num ==110 && local_vf_active==1) `toggle_tready(110)   
              else if (local_pf_num==0 && local_vf_num ==111 && local_vf_active==1) `toggle_tready(111)   
              else if (local_pf_num==0 && local_vf_num ==112 && local_vf_active==1) `toggle_tready(112)   
              else if (local_pf_num==0 && local_vf_num ==113 && local_vf_active==1) `toggle_tready(113)   
              else if (local_pf_num==0 && local_vf_num ==114 && local_vf_active==1) `toggle_tready(114)   
              else if (local_pf_num==0 && local_vf_num ==115 && local_vf_active==1) `toggle_tready(115)   
              else if (local_pf_num==0 && local_vf_num ==116 && local_vf_active==1) `toggle_tready(116)   
              else if (local_pf_num==0 && local_vf_num ==117 && local_vf_active==1) `toggle_tready(117)   
              else if (local_pf_num==0 && local_vf_num ==118 && local_vf_active==1) `toggle_tready(118)   
              else if (local_pf_num==0 && local_vf_num ==119 && local_vf_active==1) `toggle_tready(119)   
              else if (local_pf_num==0 && local_vf_num ==120 && local_vf_active==1) `toggle_tready(120)   
              else if (local_pf_num==0 && local_vf_num ==121 && local_vf_active==1) `toggle_tready(121)   
              else if (local_pf_num==0 && local_vf_num ==122 && local_vf_active==1) `toggle_tready(122)   
              else if (local_pf_num==0 && local_vf_num ==123 && local_vf_active==1) `toggle_tready(123)   
              else if (local_pf_num==0 && local_vf_num ==124 && local_vf_active==1) `toggle_tready(124)   
              else if (local_pf_num==0 && local_vf_num ==125 && local_vf_active==1) `toggle_tready(125)   
              else if (local_pf_num==0 && local_vf_num ==126 && local_vf_active==1) `toggle_tready(126)   
              else if (local_pf_num==0 && local_vf_num ==127 && local_vf_active==1) `toggle_tready(127)   
              else if (local_pf_num==0 && local_vf_num ==128 && local_vf_active==1) `toggle_tready(128)   
              else if (local_pf_num==0 && local_vf_num ==129 && local_vf_active==1) `toggle_tready(129)   
              else if (local_pf_num==0 && local_vf_num ==130 && local_vf_active==1) `toggle_tready(130)   
              else if (local_pf_num==0 && local_vf_num ==131 && local_vf_active==1) `toggle_tready(131)   
              else if (local_pf_num==0 && local_vf_num ==132 && local_vf_active==1) `toggle_tready(132)   
              else if (local_pf_num==0 && local_vf_num ==133 && local_vf_active==1) `toggle_tready(133)   
              else if (local_pf_num==0 && local_vf_num ==134 && local_vf_active==1) `toggle_tready(134)   
              else if (local_pf_num==0 && local_vf_num ==135 && local_vf_active==1) `toggle_tready(135)   
              else if (local_pf_num==0 && local_vf_num ==136 && local_vf_active==1) `toggle_tready(136)   
              else if (local_pf_num==0 && local_vf_num ==137 && local_vf_active==1) `toggle_tready(137)   
              else if (local_pf_num==0 && local_vf_num ==138 && local_vf_active==1) `toggle_tready(138)   
              else if (local_pf_num==0 && local_vf_num ==139 && local_vf_active==1) `toggle_tready(139)   
              else if (local_pf_num==0 && local_vf_num ==140 && local_vf_active==1) `toggle_tready(140)   
              else if (local_pf_num==0 && local_vf_num ==141 && local_vf_active==1) `toggle_tready(141)   
              else if (local_pf_num==0 && local_vf_num ==142 && local_vf_active==1) `toggle_tready(142)   
              else if (local_pf_num==0 && local_vf_num ==143 && local_vf_active==1) `toggle_tready(143)   
              else if (local_pf_num==0 && local_vf_num ==144 && local_vf_active==1) `toggle_tready(144)   
              else if (local_pf_num==0 && local_vf_num ==145 && local_vf_active==1) `toggle_tready(145)   
              else if (local_pf_num==0 && local_vf_num ==146 && local_vf_active==1) `toggle_tready(146)   
              else if (local_pf_num==0 && local_vf_num ==147 && local_vf_active==1) `toggle_tready(147)   
              else if (local_pf_num==0 && local_vf_num ==148 && local_vf_active==1) `toggle_tready(148)   
              else if (local_pf_num==0 && local_vf_num ==149 && local_vf_active==1) `toggle_tready(149)   
              else if (local_pf_num==0 && local_vf_num ==150 && local_vf_active==1) `toggle_tready(150)   
              else if (local_pf_num==0 && local_vf_num ==151 && local_vf_active==1) `toggle_tready(151)   
              else if (local_pf_num==0 && local_vf_num ==152 && local_vf_active==1) `toggle_tready(152)   
              else if (local_pf_num==0 && local_vf_num ==153 && local_vf_active==1) `toggle_tready(153)   
              else if (local_pf_num==0 && local_vf_num ==154 && local_vf_active==1) `toggle_tready(154)   
              else if (local_pf_num==0 && local_vf_num ==155 && local_vf_active==1) `toggle_tready(155)   
              else if (local_pf_num==0 && local_vf_num ==156 && local_vf_active==1) `toggle_tready(156)   
              else if (local_pf_num==0 && local_vf_num ==157 && local_vf_active==1) `toggle_tready(157)   
              else if (local_pf_num==0 && local_vf_num ==158 && local_vf_active==1) `toggle_tready(158)   
              else if (local_pf_num==0 && local_vf_num ==159 && local_vf_active==1) `toggle_tready(159)   
              else if (local_pf_num==0 && local_vf_num ==160 && local_vf_active==1) `toggle_tready(160)   
              else if (local_pf_num==0 && local_vf_num ==161 && local_vf_active==1) `toggle_tready(161)   
              else if (local_pf_num==0 && local_vf_num ==162 && local_vf_active==1) `toggle_tready(162)   
              else if (local_pf_num==0 && local_vf_num ==163 && local_vf_active==1) `toggle_tready(163)   
              else if (local_pf_num==0 && local_vf_num ==164 && local_vf_active==1) `toggle_tready(164)   
              else if (local_pf_num==0 && local_vf_num ==165 && local_vf_active==1) `toggle_tready(165)   
              else if (local_pf_num==0 && local_vf_num ==166 && local_vf_active==1) `toggle_tready(166)   
              else if (local_pf_num==0 && local_vf_num ==167 && local_vf_active==1) `toggle_tready(167)   
              else if (local_pf_num==0 && local_vf_num ==168 && local_vf_active==1) `toggle_tready(168)   
              else if (local_pf_num==0 && local_vf_num ==169 && local_vf_active==1) `toggle_tready(169)   
              else if (local_pf_num==0 && local_vf_num ==170 && local_vf_active==1) `toggle_tready(170)   
              else if (local_pf_num==0 && local_vf_num ==171 && local_vf_active==1) `toggle_tready(171)   
              else if (local_pf_num==0 && local_vf_num ==172 && local_vf_active==1) `toggle_tready(172)   
              else if (local_pf_num==0 && local_vf_num ==173 && local_vf_active==1) `toggle_tready(173)   
              else if (local_pf_num==0 && local_vf_num ==174 && local_vf_active==1) `toggle_tready(174)   
              else if (local_pf_num==0 && local_vf_num ==175 && local_vf_active==1) `toggle_tready(175)   
              else if (local_pf_num==0 && local_vf_num ==176 && local_vf_active==1) `toggle_tready(176)   
              else if (local_pf_num==0 && local_vf_num ==177 && local_vf_active==1) `toggle_tready(177)   
              else if (local_pf_num==0 && local_vf_num ==178 && local_vf_active==1) `toggle_tready(178)   
              else if (local_pf_num==0 && local_vf_num ==179 && local_vf_active==1) `toggle_tready(179)   
              else if (local_pf_num==0 && local_vf_num ==180 && local_vf_active==1) `toggle_tready(180)   
              else if (local_pf_num==0 && local_vf_num ==181 && local_vf_active==1) `toggle_tready(181)   
              else if (local_pf_num==0 && local_vf_num ==182 && local_vf_active==1) `toggle_tready(182)   
              else if (local_pf_num==0 && local_vf_num ==183 && local_vf_active==1) `toggle_tready(183)   
              else if (local_pf_num==0 && local_vf_num ==184 && local_vf_active==1) `toggle_tready(184)   
              else if (local_pf_num==0 && local_vf_num ==185 && local_vf_active==1) `toggle_tready(185)   
              else if (local_pf_num==0 && local_vf_num ==186 && local_vf_active==1) `toggle_tready(186)   
              else if (local_pf_num==0 && local_vf_num ==187 && local_vf_active==1) `toggle_tready(187)   
              else if (local_pf_num==0 && local_vf_num ==188 && local_vf_active==1) `toggle_tready(188)   
              else if (local_pf_num==0 && local_vf_num ==189 && local_vf_active==1) `toggle_tready(189)   
              else if (local_pf_num==0 && local_vf_num ==190 && local_vf_active==1) `toggle_tready(190)   
              else if (local_pf_num==0 && local_vf_num ==191 && local_vf_active==1) `toggle_tready(191)   
              else if (local_pf_num==0 && local_vf_num ==192 && local_vf_active==1) `toggle_tready(192)   
              else if (local_pf_num==0 && local_vf_num ==193 && local_vf_active==1) `toggle_tready(193)   
              else if (local_pf_num==0 && local_vf_num ==194 && local_vf_active==1) `toggle_tready(194)   
              else if (local_pf_num==0 && local_vf_num ==195 && local_vf_active==1) `toggle_tready(195)   
              else if (local_pf_num==0 && local_vf_num ==196 && local_vf_active==1) `toggle_tready(196)   
              else if (local_pf_num==0 && local_vf_num ==197 && local_vf_active==1) `toggle_tready(197)   
              else if (local_pf_num==0 && local_vf_num ==198 && local_vf_active==1) `toggle_tready(198)   
              else if (local_pf_num==0 && local_vf_num ==199 && local_vf_active==1) `toggle_tready(199)   
              else if (local_pf_num==0 && local_vf_num ==200 && local_vf_active==1) `toggle_tready(200)   
              else if (local_pf_num==0 && local_vf_num ==201 && local_vf_active==1) `toggle_tready(201)   
              else if (local_pf_num==0 && local_vf_num ==202 && local_vf_active==1) `toggle_tready(202)   
              else if (local_pf_num==0 && local_vf_num ==203 && local_vf_active==1) `toggle_tready(203)   
              else if (local_pf_num==0 && local_vf_num ==204 && local_vf_active==1) `toggle_tready(204)   
              else if (local_pf_num==0 && local_vf_num ==205 && local_vf_active==1) `toggle_tready(205)   
              else if (local_pf_num==0 && local_vf_num ==206 && local_vf_active==1) `toggle_tready(206)   
              else if (local_pf_num==0 && local_vf_num ==207 && local_vf_active==1) `toggle_tready(207)   
              else if (local_pf_num==0 && local_vf_num ==208 && local_vf_active==1) `toggle_tready(208)   
              else if (local_pf_num==0 && local_vf_num ==209 && local_vf_active==1) `toggle_tready(209)   
              else if (local_pf_num==0 && local_vf_num ==210 && local_vf_active==1) `toggle_tready(210)   
              else if (local_pf_num==0 && local_vf_num ==211 && local_vf_active==1) `toggle_tready(211)   
              else if (local_pf_num==0 && local_vf_num ==212 && local_vf_active==1) `toggle_tready(212)   
              else if (local_pf_num==0 && local_vf_num ==213 && local_vf_active==1) `toggle_tready(213)   
              else if (local_pf_num==0 && local_vf_num ==214 && local_vf_active==1) `toggle_tready(214)   
              else if (local_pf_num==0 && local_vf_num ==215 && local_vf_active==1) `toggle_tready(215)   
              else if (local_pf_num==0 && local_vf_num ==216 && local_vf_active==1) `toggle_tready(216)   
              else if (local_pf_num==0 && local_vf_num ==217 && local_vf_active==1) `toggle_tready(217)   
              else if (local_pf_num==0 && local_vf_num ==218 && local_vf_active==1) `toggle_tready(218)   
              else if (local_pf_num==0 && local_vf_num ==219 && local_vf_active==1) `toggle_tready(219)   
              else if (local_pf_num==0 && local_vf_num ==220 && local_vf_active==1) `toggle_tready(220)   
              else if (local_pf_num==0 && local_vf_num ==221 && local_vf_active==1) `toggle_tready(221)   
              else if (local_pf_num==0 && local_vf_num ==222 && local_vf_active==1) `toggle_tready(222)   
              else if (local_pf_num==0 && local_vf_num ==223 && local_vf_active==1) `toggle_tready(223)   
              else if (local_pf_num==0 && local_vf_num ==224 && local_vf_active==1) `toggle_tready(224)   
              else if (local_pf_num==0 && local_vf_num ==225 && local_vf_active==1) `toggle_tready(225)   
              else if (local_pf_num==0 && local_vf_num ==226 && local_vf_active==1) `toggle_tready(226)   
              else if (local_pf_num==0 && local_vf_num ==227 && local_vf_active==1) `toggle_tready(227)   
              else if (local_pf_num==0 && local_vf_num ==228 && local_vf_active==1) `toggle_tready(228)   
              else if (local_pf_num==0 && local_vf_num ==229 && local_vf_active==1) `toggle_tready(229)   
              else if (local_pf_num==0 && local_vf_num ==230 && local_vf_active==1) `toggle_tready(230)   
              else if (local_pf_num==0 && local_vf_num ==231 && local_vf_active==1) `toggle_tready(231)   
              else if (local_pf_num==0 && local_vf_num ==232 && local_vf_active==1) `toggle_tready(232)   
              else if (local_pf_num==0 && local_vf_num ==233 && local_vf_active==1) `toggle_tready(233)   
              else if (local_pf_num==0 && local_vf_num ==234 && local_vf_active==1) `toggle_tready(234)   
              else if (local_pf_num==0 && local_vf_num ==235 && local_vf_active==1) `toggle_tready(235)   
              else if (local_pf_num==0 && local_vf_num ==236 && local_vf_active==1) `toggle_tready(236)   
              else if (local_pf_num==0 && local_vf_num ==237 && local_vf_active==1) `toggle_tready(237)   
              else if (local_pf_num==0 && local_vf_num ==238 && local_vf_active==1) `toggle_tready(238)   
              else if (local_pf_num==0 && local_vf_num ==239 && local_vf_active==1) `toggle_tready(239)   
              else if (local_pf_num==0 && local_vf_num ==240 && local_vf_active==1) `toggle_tready(240)   
              else if (local_pf_num==0 && local_vf_num ==241 && local_vf_active==1) `toggle_tready(241)   
              else if (local_pf_num==0 && local_vf_num ==242 && local_vf_active==1) `toggle_tready(242)   
              else if (local_pf_num==0 && local_vf_num ==243 && local_vf_active==1) `toggle_tready(243)   
              else if (local_pf_num==0 && local_vf_num ==244 && local_vf_active==1) `toggle_tready(244)   
              else if (local_pf_num==0 && local_vf_num ==245 && local_vf_active==1) `toggle_tready(245)   
              else if (local_pf_num==0 && local_vf_num ==246 && local_vf_active==1) `toggle_tready(246)   
              else if (local_pf_num==0 && local_vf_num ==247 && local_vf_active==1) `toggle_tready(247)   
              else if (local_pf_num==0 && local_vf_num ==248 && local_vf_active==1) `toggle_tready(248)   
              else if (local_pf_num==0 && local_vf_num ==249 && local_vf_active==1) `toggle_tready(249)   
              else if (local_pf_num==0 && local_vf_num ==250 && local_vf_active==1) `toggle_tready(250)   
              else if (local_pf_num==0 && local_vf_num ==251 && local_vf_active==1) `toggle_tready(251)   
              else if (local_pf_num==0 && local_vf_num ==252 && local_vf_active==1) `toggle_tready(252)   
              else if (local_pf_num==0 && local_vf_num ==253 && local_vf_active==1) `toggle_tready(253)   
              else if (local_pf_num==0 && local_vf_num ==254 && local_vf_active==1) `toggle_tready(254)   
              else if (local_pf_num==0 && local_vf_num ==255 && local_vf_active==1) `toggle_tready(255)   
              else if (local_pf_num==0 && local_vf_num ==256 && local_vf_active==1) `toggle_tready(256)   
              else if (local_pf_num==0 && local_vf_num ==257 && local_vf_active==1) `toggle_tready(257)   
              else if (local_pf_num==0 && local_vf_num ==258 && local_vf_active==1) `toggle_tready(258)   
              else if (local_pf_num==0 && local_vf_num ==259 && local_vf_active==1) `toggle_tready(259)   
              else if (local_pf_num==0 && local_vf_num ==260 && local_vf_active==1) `toggle_tready(260)   
              else if (local_pf_num==0 && local_vf_num ==261 && local_vf_active==1) `toggle_tready(261)   
              else if (local_pf_num==0 && local_vf_num ==262 && local_vf_active==1) `toggle_tready(262)   
              else if (local_pf_num==0 && local_vf_num ==263 && local_vf_active==1) `toggle_tready(263)   
              else if (local_pf_num==0 && local_vf_num ==264 && local_vf_active==1) `toggle_tready(264)   
              else if (local_pf_num==0 && local_vf_num ==265 && local_vf_active==1) `toggle_tready(265)   
              else if (local_pf_num==0 && local_vf_num ==266 && local_vf_active==1) `toggle_tready(266)   
              else if (local_pf_num==0 && local_vf_num ==267 && local_vf_active==1) `toggle_tready(267)   
              else if (local_pf_num==0 && local_vf_num ==268 && local_vf_active==1) `toggle_tready(268)   
              else if (local_pf_num==0 && local_vf_num ==269 && local_vf_active==1) `toggle_tready(269)   
              else if (local_pf_num==0 && local_vf_num ==270 && local_vf_active==1) `toggle_tready(270)   
              else if (local_pf_num==0 && local_vf_num ==271 && local_vf_active==1) `toggle_tready(271)   
              else if (local_pf_num==0 && local_vf_num ==272 && local_vf_active==1) `toggle_tready(272)   
              else if (local_pf_num==0 && local_vf_num ==273 && local_vf_active==1) `toggle_tready(273)   
              else if (local_pf_num==0 && local_vf_num ==274 && local_vf_active==1) `toggle_tready(274)   
              else if (local_pf_num==0 && local_vf_num ==275 && local_vf_active==1) `toggle_tready(275)   
              else if (local_pf_num==0 && local_vf_num ==276 && local_vf_active==1) `toggle_tready(276)   
              else if (local_pf_num==0 && local_vf_num ==277 && local_vf_active==1) `toggle_tready(277)   
              else if (local_pf_num==0 && local_vf_num ==278 && local_vf_active==1) `toggle_tready(278)   
              else if (local_pf_num==0 && local_vf_num ==279 && local_vf_active==1) `toggle_tready(279)   
              else if (local_pf_num==0 && local_vf_num ==280 && local_vf_active==1) `toggle_tready(280)   
              else if (local_pf_num==0 && local_vf_num ==281 && local_vf_active==1) `toggle_tready(281)   
              else if (local_pf_num==0 && local_vf_num ==282 && local_vf_active==1) `toggle_tready(282)   
              else if (local_pf_num==0 && local_vf_num ==283 && local_vf_active==1) `toggle_tready(283)   
              else if (local_pf_num==0 && local_vf_num ==284 && local_vf_active==1) `toggle_tready(284)   
              else if (local_pf_num==0 && local_vf_num ==285 && local_vf_active==1) `toggle_tready(285)   
              else if (local_pf_num==0 && local_vf_num ==286 && local_vf_active==1) `toggle_tready(286)   
              else if (local_pf_num==0 && local_vf_num ==287 && local_vf_active==1) `toggle_tready(287)   
              else if (local_pf_num==0 && local_vf_num ==288 && local_vf_active==1) `toggle_tready(288)   
              else if (local_pf_num==0 && local_vf_num ==289 && local_vf_active==1) `toggle_tready(289)   
              else if (local_pf_num==0 && local_vf_num ==290 && local_vf_active==1) `toggle_tready(290)   
              else if (local_pf_num==0 && local_vf_num ==291 && local_vf_active==1) `toggle_tready(291)   
              else if (local_pf_num==0 && local_vf_num ==292 && local_vf_active==1) `toggle_tready(292)   
              else if (local_pf_num==0 && local_vf_num ==293 && local_vf_active==1) `toggle_tready(293)   
              else if (local_pf_num==0 && local_vf_num ==294 && local_vf_active==1) `toggle_tready(294)   
              else if (local_pf_num==0 && local_vf_num ==295 && local_vf_active==1) `toggle_tready(295)   
              else if (local_pf_num==0 && local_vf_num ==296 && local_vf_active==1) `toggle_tready(296)   
              else if (local_pf_num==0 && local_vf_num ==297 && local_vf_active==1) `toggle_tready(297)   
              else if (local_pf_num==0 && local_vf_num ==298 && local_vf_active==1) `toggle_tready(298)   
              else if (local_pf_num==0 && local_vf_num ==299 && local_vf_active==1) `toggle_tready(299)   
              else if (local_pf_num==0 && local_vf_num ==300 && local_vf_active==1) `toggle_tready(300)   
              else if (local_pf_num==0 && local_vf_num ==301 && local_vf_active==1) `toggle_tready(301)   
              else if (local_pf_num==0 && local_vf_num ==302 && local_vf_active==1) `toggle_tready(302)   
              else if (local_pf_num==0 && local_vf_num ==303 && local_vf_active==1) `toggle_tready(303)   
              else if (local_pf_num==0 && local_vf_num ==304 && local_vf_active==1) `toggle_tready(304)   
              else if (local_pf_num==0 && local_vf_num ==305 && local_vf_active==1) `toggle_tready(305)   
              else if (local_pf_num==0 && local_vf_num ==306 && local_vf_active==1) `toggle_tready(306)   
              else if (local_pf_num==0 && local_vf_num ==307 && local_vf_active==1) `toggle_tready(307)   
              else if (local_pf_num==0 && local_vf_num ==308 && local_vf_active==1) `toggle_tready(308)   
              else if (local_pf_num==0 && local_vf_num ==309 && local_vf_active==1) `toggle_tready(309)   
              else if (local_pf_num==0 && local_vf_num ==310 && local_vf_active==1) `toggle_tready(310)   
              else if (local_pf_num==0 && local_vf_num ==311 && local_vf_active==1) `toggle_tready(311)   
              else if (local_pf_num==0 && local_vf_num ==312 && local_vf_active==1) `toggle_tready(312)   
              else if (local_pf_num==0 && local_vf_num ==313 && local_vf_active==1) `toggle_tready(313)   
              else if (local_pf_num==0 && local_vf_num ==314 && local_vf_active==1) `toggle_tready(314)   
              else if (local_pf_num==0 && local_vf_num ==315 && local_vf_active==1) `toggle_tready(315)   
              else if (local_pf_num==0 && local_vf_num ==316 && local_vf_active==1) `toggle_tready(316)   
              else if (local_pf_num==0 && local_vf_num ==317 && local_vf_active==1) `toggle_tready(317)   
              else if (local_pf_num==0 && local_vf_num ==318 && local_vf_active==1) `toggle_tready(318)   
              else if (local_pf_num==0 && local_vf_num ==319 && local_vf_active==1) `toggle_tready(319)   
              else if (local_pf_num==0 && local_vf_num ==320 && local_vf_active==1) `toggle_tready(320)   
              else if (local_pf_num==0 && local_vf_num ==321 && local_vf_active==1) `toggle_tready(321)   
              else if (local_pf_num==0 && local_vf_num ==322 && local_vf_active==1) `toggle_tready(322)   
              else if (local_pf_num==0 && local_vf_num ==323 && local_vf_active==1) `toggle_tready(323)   
              else if (local_pf_num==0 && local_vf_num ==324 && local_vf_active==1) `toggle_tready(324)   
              else if (local_pf_num==0 && local_vf_num ==325 && local_vf_active==1) `toggle_tready(325)   
              else if (local_pf_num==0 && local_vf_num ==326 && local_vf_active==1) `toggle_tready(326)   
              else if (local_pf_num==0 && local_vf_num ==327 && local_vf_active==1) `toggle_tready(327)   
              else if (local_pf_num==0 && local_vf_num ==328 && local_vf_active==1) `toggle_tready(328)   
              else if (local_pf_num==0 && local_vf_num ==329 && local_vf_active==1) `toggle_tready(329)   
              else if (local_pf_num==0 && local_vf_num ==330 && local_vf_active==1) `toggle_tready(330)   
              else if (local_pf_num==0 && local_vf_num ==331 && local_vf_active==1) `toggle_tready(331)   
              else if (local_pf_num==0 && local_vf_num ==332 && local_vf_active==1) `toggle_tready(332)   
              else if (local_pf_num==0 && local_vf_num ==333 && local_vf_active==1) `toggle_tready(333)   
              else if (local_pf_num==0 && local_vf_num ==334 && local_vf_active==1) `toggle_tready(334)   
              else if (local_pf_num==0 && local_vf_num ==335 && local_vf_active==1) `toggle_tready(335)   
              else if (local_pf_num==0 && local_vf_num ==336 && local_vf_active==1) `toggle_tready(336)   
              else if (local_pf_num==0 && local_vf_num ==337 && local_vf_active==1) `toggle_tready(337)   
              else if (local_pf_num==0 && local_vf_num ==338 && local_vf_active==1) `toggle_tready(338)   
              else if (local_pf_num==0 && local_vf_num ==339 && local_vf_active==1) `toggle_tready(339)   
              else if (local_pf_num==0 && local_vf_num ==340 && local_vf_active==1) `toggle_tready(340)   
              else if (local_pf_num==0 && local_vf_num ==341 && local_vf_active==1) `toggle_tready(341)   
              else if (local_pf_num==0 && local_vf_num ==342 && local_vf_active==1) `toggle_tready(342)   
              else if (local_pf_num==0 && local_vf_num ==343 && local_vf_active==1) `toggle_tready(343)   
              else if (local_pf_num==0 && local_vf_num ==344 && local_vf_active==1) `toggle_tready(344)   
              else if (local_pf_num==0 && local_vf_num ==345 && local_vf_active==1) `toggle_tready(345)   
              else if (local_pf_num==0 && local_vf_num ==346 && local_vf_active==1) `toggle_tready(346)   
              else if (local_pf_num==0 && local_vf_num ==347 && local_vf_active==1) `toggle_tready(347)   
              else if (local_pf_num==0 && local_vf_num ==348 && local_vf_active==1) `toggle_tready(348)   
              else if (local_pf_num==0 && local_vf_num ==349 && local_vf_active==1) `toggle_tready(349)   
              else if (local_pf_num==0 && local_vf_num ==350 && local_vf_active==1) `toggle_tready(350)   
              else if (local_pf_num==0 && local_vf_num ==351 && local_vf_active==1) `toggle_tready(351)   
              else if (local_pf_num==0 && local_vf_num ==352 && local_vf_active==1) `toggle_tready(352)   
              else if (local_pf_num==0 && local_vf_num ==353 && local_vf_active==1) `toggle_tready(353)   
              else if (local_pf_num==0 && local_vf_num ==354 && local_vf_active==1) `toggle_tready(354)   
              else if (local_pf_num==0 && local_vf_num ==355 && local_vf_active==1) `toggle_tready(355)   
              else if (local_pf_num==0 && local_vf_num ==356 && local_vf_active==1) `toggle_tready(356)   
              else if (local_pf_num==0 && local_vf_num ==357 && local_vf_active==1) `toggle_tready(357)   
              else if (local_pf_num==0 && local_vf_num ==358 && local_vf_active==1) `toggle_tready(358)   
              else if (local_pf_num==0 && local_vf_num ==359 && local_vf_active==1) `toggle_tready(359)   
              else if (local_pf_num==0 && local_vf_num ==360 && local_vf_active==1) `toggle_tready(360)   
              else if (local_pf_num==0 && local_vf_num ==361 && local_vf_active==1) `toggle_tready(361)   
              else if (local_pf_num==0 && local_vf_num ==362 && local_vf_active==1) `toggle_tready(362)   
              else if (local_pf_num==0 && local_vf_num ==363 && local_vf_active==1) `toggle_tready(363)   
              else if (local_pf_num==0 && local_vf_num ==364 && local_vf_active==1) `toggle_tready(364)   
              else if (local_pf_num==0 && local_vf_num ==365 && local_vf_active==1) `toggle_tready(365)   
              else if (local_pf_num==0 && local_vf_num ==366 && local_vf_active==1) `toggle_tready(366)   
              else if (local_pf_num==0 && local_vf_num ==367 && local_vf_active==1) `toggle_tready(367)   
              else if (local_pf_num==0 && local_vf_num ==368 && local_vf_active==1) `toggle_tready(368)   
              else if (local_pf_num==0 && local_vf_num ==369 && local_vf_active==1) `toggle_tready(369)   
              else if (local_pf_num==0 && local_vf_num ==370 && local_vf_active==1) `toggle_tready(370)   
              else if (local_pf_num==0 && local_vf_num ==371 && local_vf_active==1) `toggle_tready(371)   
              else if (local_pf_num==0 && local_vf_num ==372 && local_vf_active==1) `toggle_tready(372)   
              else if (local_pf_num==0 && local_vf_num ==373 && local_vf_active==1) `toggle_tready(373)   
              else if (local_pf_num==0 && local_vf_num ==374 && local_vf_active==1) `toggle_tready(374)   
              else if (local_pf_num==0 && local_vf_num ==375 && local_vf_active==1) `toggle_tready(375)   
              else if (local_pf_num==0 && local_vf_num ==376 && local_vf_active==1) `toggle_tready(376)   
              else if (local_pf_num==0 && local_vf_num ==377 && local_vf_active==1) `toggle_tready(377)   
              else if (local_pf_num==0 && local_vf_num ==378 && local_vf_active==1) `toggle_tready(378)   
              else if (local_pf_num==0 && local_vf_num ==379 && local_vf_active==1) `toggle_tready(379)   
              else if (local_pf_num==0 && local_vf_num ==380 && local_vf_active==1) `toggle_tready(380)   
              else if (local_pf_num==0 && local_vf_num ==381 && local_vf_active==1) `toggle_tready(381)   
              else if (local_pf_num==0 && local_vf_num ==382 && local_vf_active==1) `toggle_tready(382)   
              else if (local_pf_num==0 && local_vf_num ==383 && local_vf_active==1) `toggle_tready(383)   
              else if (local_pf_num==0 && local_vf_num ==384 && local_vf_active==1) `toggle_tready(384)   
              else if (local_pf_num==0 && local_vf_num ==385 && local_vf_active==1) `toggle_tready(385)   
              else if (local_pf_num==0 && local_vf_num ==386 && local_vf_active==1) `toggle_tready(386)   
              else if (local_pf_num==0 && local_vf_num ==387 && local_vf_active==1) `toggle_tready(387)   
              else if (local_pf_num==0 && local_vf_num ==388 && local_vf_active==1) `toggle_tready(388)   
              else if (local_pf_num==0 && local_vf_num ==389 && local_vf_active==1) `toggle_tready(389)   
              else if (local_pf_num==0 && local_vf_num ==390 && local_vf_active==1) `toggle_tready(390)   
              else if (local_pf_num==0 && local_vf_num ==391 && local_vf_active==1) `toggle_tready(391)   
              else if (local_pf_num==0 && local_vf_num ==392 && local_vf_active==1) `toggle_tready(392)   
              else if (local_pf_num==0 && local_vf_num ==393 && local_vf_active==1) `toggle_tready(393)   
              else if (local_pf_num==0 && local_vf_num ==394 && local_vf_active==1) `toggle_tready(394)   
              else if (local_pf_num==0 && local_vf_num ==395 && local_vf_active==1) `toggle_tready(395)   
              else if (local_pf_num==0 && local_vf_num ==396 && local_vf_active==1) `toggle_tready(396)   
              else if (local_pf_num==0 && local_vf_num ==397 && local_vf_active==1) `toggle_tready(397)   
              else if (local_pf_num==0 && local_vf_num ==398 && local_vf_active==1) `toggle_tready(398)   
              else if (local_pf_num==0 && local_vf_num ==399 && local_vf_active==1) `toggle_tready(399)   
              else if (local_pf_num==0 && local_vf_num ==400 && local_vf_active==1) `toggle_tready(400)   
              else if (local_pf_num==0 && local_vf_num ==401 && local_vf_active==1) `toggle_tready(401)   
              else if (local_pf_num==0 && local_vf_num ==402 && local_vf_active==1) `toggle_tready(402)   
              else if (local_pf_num==0 && local_vf_num ==403 && local_vf_active==1) `toggle_tready(403)   
              else if (local_pf_num==0 && local_vf_num ==404 && local_vf_active==1) `toggle_tready(404)   
              else if (local_pf_num==0 && local_vf_num ==405 && local_vf_active==1) `toggle_tready(405)   
              else if (local_pf_num==0 && local_vf_num ==406 && local_vf_active==1) `toggle_tready(406)   
              else if (local_pf_num==0 && local_vf_num ==407 && local_vf_active==1) `toggle_tready(407)   
              else if (local_pf_num==0 && local_vf_num ==408 && local_vf_active==1) `toggle_tready(408)   
              else if (local_pf_num==0 && local_vf_num ==409 && local_vf_active==1) `toggle_tready(409)   
              else if (local_pf_num==0 && local_vf_num ==410 && local_vf_active==1) `toggle_tready(410)   
              else if (local_pf_num==0 && local_vf_num ==411 && local_vf_active==1) `toggle_tready(411)   
              else if (local_pf_num==0 && local_vf_num ==412 && local_vf_active==1) `toggle_tready(412)   
              else if (local_pf_num==0 && local_vf_num ==413 && local_vf_active==1) `toggle_tready(413)   
              else if (local_pf_num==0 && local_vf_num ==414 && local_vf_active==1) `toggle_tready(414)   
              else if (local_pf_num==0 && local_vf_num ==415 && local_vf_active==1) `toggle_tready(415)   
              else if (local_pf_num==0 && local_vf_num ==416 && local_vf_active==1) `toggle_tready(416)   
              else if (local_pf_num==0 && local_vf_num ==417 && local_vf_active==1) `toggle_tready(417)   
              else if (local_pf_num==0 && local_vf_num ==418 && local_vf_active==1) `toggle_tready(418)   
              else if (local_pf_num==0 && local_vf_num ==419 && local_vf_active==1) `toggle_tready(419)   
              else if (local_pf_num==0 && local_vf_num ==420 && local_vf_active==1) `toggle_tready(420)   
              else if (local_pf_num==0 && local_vf_num ==421 && local_vf_active==1) `toggle_tready(421)   
              else if (local_pf_num==0 && local_vf_num ==422 && local_vf_active==1) `toggle_tready(422)   
              else if (local_pf_num==0 && local_vf_num ==423 && local_vf_active==1) `toggle_tready(423)   
              else if (local_pf_num==0 && local_vf_num ==424 && local_vf_active==1) `toggle_tready(424)   
              else if (local_pf_num==0 && local_vf_num ==425 && local_vf_active==1) `toggle_tready(425)   
              else if (local_pf_num==0 && local_vf_num ==426 && local_vf_active==1) `toggle_tready(426)   
              else if (local_pf_num==0 && local_vf_num ==427 && local_vf_active==1) `toggle_tready(427)   
              else if (local_pf_num==0 && local_vf_num ==428 && local_vf_active==1) `toggle_tready(428)   
              else if (local_pf_num==0 && local_vf_num ==429 && local_vf_active==1) `toggle_tready(429)   
              else if (local_pf_num==0 && local_vf_num ==430 && local_vf_active==1) `toggle_tready(430)   
              else if (local_pf_num==0 && local_vf_num ==431 && local_vf_active==1) `toggle_tready(431)   
              else if (local_pf_num==0 && local_vf_num ==432 && local_vf_active==1) `toggle_tready(432)   
              else if (local_pf_num==0 && local_vf_num ==433 && local_vf_active==1) `toggle_tready(433)   
              else if (local_pf_num==0 && local_vf_num ==434 && local_vf_active==1) `toggle_tready(434)   
              else if (local_pf_num==0 && local_vf_num ==435 && local_vf_active==1) `toggle_tready(435)   
              else if (local_pf_num==0 && local_vf_num ==436 && local_vf_active==1) `toggle_tready(436)   
              else if (local_pf_num==0 && local_vf_num ==437 && local_vf_active==1) `toggle_tready(437)   
              else if (local_pf_num==0 && local_vf_num ==438 && local_vf_active==1) `toggle_tready(438)   
              else if (local_pf_num==0 && local_vf_num ==439 && local_vf_active==1) `toggle_tready(439)   
              else if (local_pf_num==0 && local_vf_num ==440 && local_vf_active==1) `toggle_tready(440)   
              else if (local_pf_num==0 && local_vf_num ==441 && local_vf_active==1) `toggle_tready(441)   
              else if (local_pf_num==0 && local_vf_num ==442 && local_vf_active==1) `toggle_tready(442)   
              else if (local_pf_num==0 && local_vf_num ==443 && local_vf_active==1) `toggle_tready(443)   
              else if (local_pf_num==0 && local_vf_num ==444 && local_vf_active==1) `toggle_tready(444)   
              else if (local_pf_num==0 && local_vf_num ==445 && local_vf_active==1) `toggle_tready(445)   
              else if (local_pf_num==0 && local_vf_num ==446 && local_vf_active==1) `toggle_tready(446)   
              else if (local_pf_num==0 && local_vf_num ==447 && local_vf_active==1) `toggle_tready(447)   
              else if (local_pf_num==0 && local_vf_num ==448 && local_vf_active==1) `toggle_tready(448)   
              else if (local_pf_num==0 && local_vf_num ==449 && local_vf_active==1) `toggle_tready(449)   
              else if (local_pf_num==0 && local_vf_num ==450 && local_vf_active==1) `toggle_tready(450)   
              else if (local_pf_num==0 && local_vf_num ==451 && local_vf_active==1) `toggle_tready(451)   
              else if (local_pf_num==0 && local_vf_num ==452 && local_vf_active==1) `toggle_tready(452)   
              else if (local_pf_num==0 && local_vf_num ==453 && local_vf_active==1) `toggle_tready(453)   
              else if (local_pf_num==0 && local_vf_num ==454 && local_vf_active==1) `toggle_tready(454)   
              else if (local_pf_num==0 && local_vf_num ==455 && local_vf_active==1) `toggle_tready(455)   
              else if (local_pf_num==0 && local_vf_num ==456 && local_vf_active==1) `toggle_tready(456)   
              else if (local_pf_num==0 && local_vf_num ==457 && local_vf_active==1) `toggle_tready(457)   
              else if (local_pf_num==0 && local_vf_num ==458 && local_vf_active==1) `toggle_tready(458)   
              else if (local_pf_num==0 && local_vf_num ==459 && local_vf_active==1) `toggle_tready(459)   
              else if (local_pf_num==0 && local_vf_num ==460 && local_vf_active==1) `toggle_tready(460)   
              else if (local_pf_num==0 && local_vf_num ==461 && local_vf_active==1) `toggle_tready(461)   
              else if (local_pf_num==0 && local_vf_num ==462 && local_vf_active==1) `toggle_tready(462)   
              else if (local_pf_num==0 && local_vf_num ==463 && local_vf_active==1) `toggle_tready(463)   
              else if (local_pf_num==0 && local_vf_num ==464 && local_vf_active==1) `toggle_tready(464)   
              else if (local_pf_num==0 && local_vf_num ==465 && local_vf_active==1) `toggle_tready(465)   
              else if (local_pf_num==0 && local_vf_num ==466 && local_vf_active==1) `toggle_tready(466)   
              else if (local_pf_num==0 && local_vf_num ==467 && local_vf_active==1) `toggle_tready(467)   
              else if (local_pf_num==0 && local_vf_num ==468 && local_vf_active==1) `toggle_tready(468)   
              else if (local_pf_num==0 && local_vf_num ==469 && local_vf_active==1) `toggle_tready(469)   
              else if (local_pf_num==0 && local_vf_num ==470 && local_vf_active==1) `toggle_tready(470)   
              else if (local_pf_num==0 && local_vf_num ==471 && local_vf_active==1) `toggle_tready(471)   
              else if (local_pf_num==0 && local_vf_num ==472 && local_vf_active==1) `toggle_tready(472)   
              else if (local_pf_num==0 && local_vf_num ==473 && local_vf_active==1) `toggle_tready(473)   
              else if (local_pf_num==0 && local_vf_num ==474 && local_vf_active==1) `toggle_tready(474)   
              else if (local_pf_num==0 && local_vf_num ==475 && local_vf_active==1) `toggle_tready(475)   
              else if (local_pf_num==0 && local_vf_num ==476 && local_vf_active==1) `toggle_tready(476)   
              else if (local_pf_num==0 && local_vf_num ==477 && local_vf_active==1) `toggle_tready(477)   
              else if (local_pf_num==0 && local_vf_num ==478 && local_vf_active==1) `toggle_tready(478)   
              else if (local_pf_num==0 && local_vf_num ==479 && local_vf_active==1) `toggle_tready(479)   
              else if (local_pf_num==0 && local_vf_num ==480 && local_vf_active==1) `toggle_tready(480)   
              else if (local_pf_num==0 && local_vf_num ==481 && local_vf_active==1) `toggle_tready(481)   
              else if (local_pf_num==0 && local_vf_num ==482 && local_vf_active==1) `toggle_tready(482)   
              else if (local_pf_num==0 && local_vf_num ==483 && local_vf_active==1) `toggle_tready(483)   
              else if (local_pf_num==0 && local_vf_num ==484 && local_vf_active==1) `toggle_tready(484)   
              else if (local_pf_num==0 && local_vf_num ==485 && local_vf_active==1) `toggle_tready(485)   
              else if (local_pf_num==0 && local_vf_num ==486 && local_vf_active==1) `toggle_tready(486)   
              else if (local_pf_num==0 && local_vf_num ==487 && local_vf_active==1) `toggle_tready(487)   
              else if (local_pf_num==0 && local_vf_num ==488 && local_vf_active==1) `toggle_tready(488)   
              else if (local_pf_num==0 && local_vf_num ==489 && local_vf_active==1) `toggle_tready(489)   
              else if (local_pf_num==0 && local_vf_num ==490 && local_vf_active==1) `toggle_tready(490)   
              else if (local_pf_num==0 && local_vf_num ==491 && local_vf_active==1) `toggle_tready(491)   
              else if (local_pf_num==0 && local_vf_num ==492 && local_vf_active==1) `toggle_tready(492)   
              else if (local_pf_num==0 && local_vf_num ==493 && local_vf_active==1) `toggle_tready(493)   
              else if (local_pf_num==0 && local_vf_num ==494 && local_vf_active==1) `toggle_tready(494)   
              else if (local_pf_num==0 && local_vf_num ==495 && local_vf_active==1) `toggle_tready(495)   
              else if (local_pf_num==0 && local_vf_num ==496 && local_vf_active==1) `toggle_tready(496)   
              else if (local_pf_num==0 && local_vf_num ==497 && local_vf_active==1) `toggle_tready(497)   
              else if (local_pf_num==0 && local_vf_num ==498 && local_vf_active==1) `toggle_tready(498)   
              else if (local_pf_num==0 && local_vf_num ==499 && local_vf_active==1) `toggle_tready(499)   
              else if (local_pf_num==0 && local_vf_num ==500 && local_vf_active==1) `toggle_tready(500)   
              else if (local_pf_num==0 && local_vf_num ==501 && local_vf_active==1) `toggle_tready(501)   
              else if (local_pf_num==0 && local_vf_num ==502 && local_vf_active==1) `toggle_tready(502)   
              else if (local_pf_num==0 && local_vf_num ==503 && local_vf_active==1) `toggle_tready(503)   
              else if (local_pf_num==0 && local_vf_num ==504 && local_vf_active==1) `toggle_tready(504)   
              else if (local_pf_num==0 && local_vf_num ==505 && local_vf_active==1) `toggle_tready(505)   
              else if (local_pf_num==0 && local_vf_num ==506 && local_vf_active==1) `toggle_tready(506)   
              else if (local_pf_num==0 && local_vf_num ==507 && local_vf_active==1) `toggle_tready(507)   
              else if (local_pf_num==0 && local_vf_num ==508 && local_vf_active==1) `toggle_tready(508)   
              else if (local_pf_num==0 && local_vf_num ==509 && local_vf_active==1) `toggle_tready(509)   
              else if (local_pf_num==0 && local_vf_num ==510 && local_vf_active==1) `toggle_tready(510)   
              else if (local_pf_num==0 && local_vf_num ==511 && local_vf_active==1) `toggle_tready(511)   
              else if (local_pf_num==0 && local_vf_num ==512 && local_vf_active==1) `toggle_tready(512)   
              else if (local_pf_num==0 && local_vf_num ==513 && local_vf_active==1) `toggle_tready(513)   
              else if (local_pf_num==0 && local_vf_num ==514 && local_vf_active==1) `toggle_tready(514)   
              else if (local_pf_num==0 && local_vf_num ==515 && local_vf_active==1) `toggle_tready(515)   
              else if (local_pf_num==0 && local_vf_num ==516 && local_vf_active==1) `toggle_tready(516)   
              else if (local_pf_num==0 && local_vf_num ==517 && local_vf_active==1) `toggle_tready(517)   
              else if (local_pf_num==0 && local_vf_num ==518 && local_vf_active==1) `toggle_tready(518)   
              else if (local_pf_num==0 && local_vf_num ==519 && local_vf_active==1) `toggle_tready(519)   
              else if (local_pf_num==0 && local_vf_num ==520 && local_vf_active==1) `toggle_tready(520)   
              else if (local_pf_num==0 && local_vf_num ==521 && local_vf_active==1) `toggle_tready(521)   
              else if (local_pf_num==0 && local_vf_num ==522 && local_vf_active==1) `toggle_tready(522)   
              else if (local_pf_num==0 && local_vf_num ==523 && local_vf_active==1) `toggle_tready(523)   
              else if (local_pf_num==0 && local_vf_num ==524 && local_vf_active==1) `toggle_tready(524)   
              else if (local_pf_num==0 && local_vf_num ==525 && local_vf_active==1) `toggle_tready(525)   
              else if (local_pf_num==0 && local_vf_num ==526 && local_vf_active==1) `toggle_tready(526)   
              else if (local_pf_num==0 && local_vf_num ==527 && local_vf_active==1) `toggle_tready(527)   
              else if (local_pf_num==0 && local_vf_num ==528 && local_vf_active==1) `toggle_tready(528)   
              else if (local_pf_num==0 && local_vf_num ==529 && local_vf_active==1) `toggle_tready(529)   
              else if (local_pf_num==0 && local_vf_num ==530 && local_vf_active==1) `toggle_tready(530)   
              else if (local_pf_num==0 && local_vf_num ==531 && local_vf_active==1) `toggle_tready(531)   
              else if (local_pf_num==0 && local_vf_num ==532 && local_vf_active==1) `toggle_tready(532)   
              else if (local_pf_num==0 && local_vf_num ==533 && local_vf_active==1) `toggle_tready(533)   
              else if (local_pf_num==0 && local_vf_num ==534 && local_vf_active==1) `toggle_tready(534)   
              else if (local_pf_num==0 && local_vf_num ==535 && local_vf_active==1) `toggle_tready(535)   
              else if (local_pf_num==0 && local_vf_num ==536 && local_vf_active==1) `toggle_tready(536)   
              else if (local_pf_num==0 && local_vf_num ==537 && local_vf_active==1) `toggle_tready(537)   
              else if (local_pf_num==0 && local_vf_num ==538 && local_vf_active==1) `toggle_tready(538)   
              else if (local_pf_num==0 && local_vf_num ==539 && local_vf_active==1) `toggle_tready(539)   
              else if (local_pf_num==0 && local_vf_num ==540 && local_vf_active==1) `toggle_tready(540)   
              else if (local_pf_num==0 && local_vf_num ==541 && local_vf_active==1) `toggle_tready(541)   
              else if (local_pf_num==0 && local_vf_num ==542 && local_vf_active==1) `toggle_tready(542)   
              else if (local_pf_num==0 && local_vf_num ==543 && local_vf_active==1) `toggle_tready(543)   
              else if (local_pf_num==0 && local_vf_num ==544 && local_vf_active==1) `toggle_tready(544)   
              else if (local_pf_num==0 && local_vf_num ==545 && local_vf_active==1) `toggle_tready(545)   
              else if (local_pf_num==0 && local_vf_num ==546 && local_vf_active==1) `toggle_tready(546)   
              else if (local_pf_num==0 && local_vf_num ==547 && local_vf_active==1) `toggle_tready(547)   
              else if (local_pf_num==0 && local_vf_num ==548 && local_vf_active==1) `toggle_tready(548)   
              else if (local_pf_num==0 && local_vf_num ==549 && local_vf_active==1) `toggle_tready(549)   
              else if (local_pf_num==0 && local_vf_num ==550 && local_vf_active==1) `toggle_tready(550)   
              else if (local_pf_num==0 && local_vf_num ==551 && local_vf_active==1) `toggle_tready(551)   
              else if (local_pf_num==0 && local_vf_num ==552 && local_vf_active==1) `toggle_tready(552)   
              else if (local_pf_num==0 && local_vf_num ==553 && local_vf_active==1) `toggle_tready(553)   
              else if (local_pf_num==0 && local_vf_num ==554 && local_vf_active==1) `toggle_tready(554)   
              else if (local_pf_num==0 && local_vf_num ==555 && local_vf_active==1) `toggle_tready(555)   
              else if (local_pf_num==0 && local_vf_num ==556 && local_vf_active==1) `toggle_tready(556)   
              else if (local_pf_num==0 && local_vf_num ==557 && local_vf_active==1) `toggle_tready(557)   
              else if (local_pf_num==0 && local_vf_num ==558 && local_vf_active==1) `toggle_tready(558)   
              else if (local_pf_num==0 && local_vf_num ==559 && local_vf_active==1) `toggle_tready(559)   
              else if (local_pf_num==0 && local_vf_num ==560 && local_vf_active==1) `toggle_tready(560)   
              else if (local_pf_num==0 && local_vf_num ==561 && local_vf_active==1) `toggle_tready(561)   
              else if (local_pf_num==0 && local_vf_num ==562 && local_vf_active==1) `toggle_tready(562)   
              else if (local_pf_num==0 && local_vf_num ==563 && local_vf_active==1) `toggle_tready(563)   
              else if (local_pf_num==0 && local_vf_num ==564 && local_vf_active==1) `toggle_tready(564)   
              else if (local_pf_num==0 && local_vf_num ==565 && local_vf_active==1) `toggle_tready(565)   
              else if (local_pf_num==0 && local_vf_num ==566 && local_vf_active==1) `toggle_tready(566)   
              else if (local_pf_num==0 && local_vf_num ==567 && local_vf_active==1) `toggle_tready(567)   
              else if (local_pf_num==0 && local_vf_num ==568 && local_vf_active==1) `toggle_tready(568)   
              else if (local_pf_num==0 && local_vf_num ==569 && local_vf_active==1) `toggle_tready(569)   
              else if (local_pf_num==0 && local_vf_num ==570 && local_vf_active==1) `toggle_tready(570)   
              else if (local_pf_num==0 && local_vf_num ==571 && local_vf_active==1) `toggle_tready(571)   
              else if (local_pf_num==0 && local_vf_num ==572 && local_vf_active==1) `toggle_tready(572)   
              else if (local_pf_num==0 && local_vf_num ==573 && local_vf_active==1) `toggle_tready(573)   
              else if (local_pf_num==0 && local_vf_num ==574 && local_vf_active==1) `toggle_tready(574)   
              else if (local_pf_num==0 && local_vf_num ==575 && local_vf_active==1) `toggle_tready(575)   
              else if (local_pf_num==0 && local_vf_num ==576 && local_vf_active==1) `toggle_tready(576)   
              else if (local_pf_num==0 && local_vf_num ==577 && local_vf_active==1) `toggle_tready(577)   
              else if (local_pf_num==0 && local_vf_num ==578 && local_vf_active==1) `toggle_tready(578)   
              else if (local_pf_num==0 && local_vf_num ==579 && local_vf_active==1) `toggle_tready(579)   
              else if (local_pf_num==0 && local_vf_num ==580 && local_vf_active==1) `toggle_tready(580)   
              else if (local_pf_num==0 && local_vf_num ==581 && local_vf_active==1) `toggle_tready(581)   
              else if (local_pf_num==0 && local_vf_num ==582 && local_vf_active==1) `toggle_tready(582)   
              else if (local_pf_num==0 && local_vf_num ==583 && local_vf_active==1) `toggle_tready(583)   
              else if (local_pf_num==0 && local_vf_num ==584 && local_vf_active==1) `toggle_tready(584)   
              else if (local_pf_num==0 && local_vf_num ==585 && local_vf_active==1) `toggle_tready(585)   
              else if (local_pf_num==0 && local_vf_num ==586 && local_vf_active==1) `toggle_tready(586)   
              else if (local_pf_num==0 && local_vf_num ==587 && local_vf_active==1) `toggle_tready(587)   
              else if (local_pf_num==0 && local_vf_num ==588 && local_vf_active==1) `toggle_tready(588)   
              else if (local_pf_num==0 && local_vf_num ==589 && local_vf_active==1) `toggle_tready(589)   
              else if (local_pf_num==0 && local_vf_num ==590 && local_vf_active==1) `toggle_tready(590)   
              else if (local_pf_num==0 && local_vf_num ==591 && local_vf_active==1) `toggle_tready(591)   
              else if (local_pf_num==0 && local_vf_num ==592 && local_vf_active==1) `toggle_tready(592)   
              else if (local_pf_num==0 && local_vf_num ==593 && local_vf_active==1) `toggle_tready(593)   
              else if (local_pf_num==0 && local_vf_num ==594 && local_vf_active==1) `toggle_tready(594)   
              else if (local_pf_num==0 && local_vf_num ==595 && local_vf_active==1) `toggle_tready(595)   
              else if (local_pf_num==0 && local_vf_num ==596 && local_vf_active==1) `toggle_tready(596)   
              else if (local_pf_num==0 && local_vf_num ==597 && local_vf_active==1) `toggle_tready(597)   
              else if (local_pf_num==0 && local_vf_num ==598 && local_vf_active==1) `toggle_tready(598)   
              else if (local_pf_num==0 && local_vf_num ==599 && local_vf_active==1) `toggle_tready(599)   
              else if (local_pf_num==0 && local_vf_num ==600 && local_vf_active==1) `toggle_tready(600)   
              else if (local_pf_num==0 && local_vf_num ==601 && local_vf_active==1) `toggle_tready(601)   
              else if (local_pf_num==0 && local_vf_num ==602 && local_vf_active==1) `toggle_tready(602)   
              else if (local_pf_num==0 && local_vf_num ==603 && local_vf_active==1) `toggle_tready(603)   
              else if (local_pf_num==0 && local_vf_num ==604 && local_vf_active==1) `toggle_tready(604)   
              else if (local_pf_num==0 && local_vf_num ==605 && local_vf_active==1) `toggle_tready(605)   
              else if (local_pf_num==0 && local_vf_num ==606 && local_vf_active==1) `toggle_tready(606)   
              else if (local_pf_num==0 && local_vf_num ==607 && local_vf_active==1) `toggle_tready(607)   
              else if (local_pf_num==0 && local_vf_num ==608 && local_vf_active==1) `toggle_tready(608)   
              else if (local_pf_num==0 && local_vf_num ==609 && local_vf_active==1) `toggle_tready(609)   
              else if (local_pf_num==0 && local_vf_num ==610 && local_vf_active==1) `toggle_tready(610)   
              else if (local_pf_num==0 && local_vf_num ==611 && local_vf_active==1) `toggle_tready(611)   
              else if (local_pf_num==0 && local_vf_num ==612 && local_vf_active==1) `toggle_tready(612)   
              else if (local_pf_num==0 && local_vf_num ==613 && local_vf_active==1) `toggle_tready(613)   
              else if (local_pf_num==0 && local_vf_num ==614 && local_vf_active==1) `toggle_tready(614)   
              else if (local_pf_num==0 && local_vf_num ==615 && local_vf_active==1) `toggle_tready(615)   
              else if (local_pf_num==0 && local_vf_num ==616 && local_vf_active==1) `toggle_tready(616)   
              else if (local_pf_num==0 && local_vf_num ==617 && local_vf_active==1) `toggle_tready(617)   
              else if (local_pf_num==0 && local_vf_num ==618 && local_vf_active==1) `toggle_tready(618)   
              else if (local_pf_num==0 && local_vf_num ==619 && local_vf_active==1) `toggle_tready(619)   
              else if (local_pf_num==0 && local_vf_num ==620 && local_vf_active==1) `toggle_tready(620)   
              else if (local_pf_num==0 && local_vf_num ==621 && local_vf_active==1) `toggle_tready(621)   
              else if (local_pf_num==0 && local_vf_num ==622 && local_vf_active==1) `toggle_tready(622)   
              else if (local_pf_num==0 && local_vf_num ==623 && local_vf_active==1) `toggle_tready(623)   
              else if (local_pf_num==0 && local_vf_num ==624 && local_vf_active==1) `toggle_tready(624)   
              else if (local_pf_num==0 && local_vf_num ==625 && local_vf_active==1) `toggle_tready(625)   
              else if (local_pf_num==0 && local_vf_num ==626 && local_vf_active==1) `toggle_tready(626)   
              else if (local_pf_num==0 && local_vf_num ==627 && local_vf_active==1) `toggle_tready(627)   
              else if (local_pf_num==0 && local_vf_num ==628 && local_vf_active==1) `toggle_tready(628)   
              else if (local_pf_num==0 && local_vf_num ==629 && local_vf_active==1) `toggle_tready(629)   
              else if (local_pf_num==0 && local_vf_num ==630 && local_vf_active==1) `toggle_tready(630)   
              else if (local_pf_num==0 && local_vf_num ==631 && local_vf_active==1) `toggle_tready(631)   
              else if (local_pf_num==0 && local_vf_num ==632 && local_vf_active==1) `toggle_tready(632)   
              else if (local_pf_num==0 && local_vf_num ==633 && local_vf_active==1) `toggle_tready(633)   
              else if (local_pf_num==0 && local_vf_num ==634 && local_vf_active==1) `toggle_tready(634)   
              else if (local_pf_num==0 && local_vf_num ==635 && local_vf_active==1) `toggle_tready(635)   
              else if (local_pf_num==0 && local_vf_num ==636 && local_vf_active==1) `toggle_tready(636)   
              else if (local_pf_num==0 && local_vf_num ==637 && local_vf_active==1) `toggle_tready(637)   
              else if (local_pf_num==0 && local_vf_num ==638 && local_vf_active==1) `toggle_tready(638)   
              else if (local_pf_num==0 && local_vf_num ==639 && local_vf_active==1) `toggle_tready(639)   
              else if (local_pf_num==0 && local_vf_num ==640 && local_vf_active==1) `toggle_tready(640)   
              else if (local_pf_num==0 && local_vf_num ==641 && local_vf_active==1) `toggle_tready(641)   
              else if (local_pf_num==0 && local_vf_num ==642 && local_vf_active==1) `toggle_tready(642)   
              else if (local_pf_num==0 && local_vf_num ==643 && local_vf_active==1) `toggle_tready(643)   
              else if (local_pf_num==0 && local_vf_num ==644 && local_vf_active==1) `toggle_tready(644)   
              else if (local_pf_num==0 && local_vf_num ==645 && local_vf_active==1) `toggle_tready(645)   
              else if (local_pf_num==0 && local_vf_num ==646 && local_vf_active==1) `toggle_tready(646)   
              else if (local_pf_num==0 && local_vf_num ==647 && local_vf_active==1) `toggle_tready(647)   
              else if (local_pf_num==0 && local_vf_num ==648 && local_vf_active==1) `toggle_tready(648)   
              else if (local_pf_num==0 && local_vf_num ==649 && local_vf_active==1) `toggle_tready(649)   
              else if (local_pf_num==0 && local_vf_num ==650 && local_vf_active==1) `toggle_tready(650)   
              else if (local_pf_num==0 && local_vf_num ==651 && local_vf_active==1) `toggle_tready(651)   
              else if (local_pf_num==0 && local_vf_num ==652 && local_vf_active==1) `toggle_tready(652)   
              else if (local_pf_num==0 && local_vf_num ==653 && local_vf_active==1) `toggle_tready(653)   
              else if (local_pf_num==0 && local_vf_num ==654 && local_vf_active==1) `toggle_tready(654)   
              else if (local_pf_num==0 && local_vf_num ==655 && local_vf_active==1) `toggle_tready(655)   
              else if (local_pf_num==0 && local_vf_num ==656 && local_vf_active==1) `toggle_tready(656)   
              else if (local_pf_num==0 && local_vf_num ==657 && local_vf_active==1) `toggle_tready(657)   
              else if (local_pf_num==0 && local_vf_num ==658 && local_vf_active==1) `toggle_tready(658)   
              else if (local_pf_num==0 && local_vf_num ==659 && local_vf_active==1) `toggle_tready(659)   
              else if (local_pf_num==0 && local_vf_num ==660 && local_vf_active==1) `toggle_tready(660)   
              else if (local_pf_num==0 && local_vf_num ==661 && local_vf_active==1) `toggle_tready(661)   
              else if (local_pf_num==0 && local_vf_num ==662 && local_vf_active==1) `toggle_tready(662)   
              else if (local_pf_num==0 && local_vf_num ==663 && local_vf_active==1) `toggle_tready(663)   
              else if (local_pf_num==0 && local_vf_num ==664 && local_vf_active==1) `toggle_tready(664)   
              else if (local_pf_num==0 && local_vf_num ==665 && local_vf_active==1) `toggle_tready(665)   
              else if (local_pf_num==0 && local_vf_num ==666 && local_vf_active==1) `toggle_tready(666)   
              else if (local_pf_num==0 && local_vf_num ==667 && local_vf_active==1) `toggle_tready(667)   
              else if (local_pf_num==0 && local_vf_num ==668 && local_vf_active==1) `toggle_tready(668)   
              else if (local_pf_num==0 && local_vf_num ==669 && local_vf_active==1) `toggle_tready(669)   
              else if (local_pf_num==0 && local_vf_num ==670 && local_vf_active==1) `toggle_tready(670)   
              else if (local_pf_num==0 && local_vf_num ==671 && local_vf_active==1) `toggle_tready(671)   
              else if (local_pf_num==0 && local_vf_num ==672 && local_vf_active==1) `toggle_tready(672)   
              else if (local_pf_num==0 && local_vf_num ==673 && local_vf_active==1) `toggle_tready(673)   
              else if (local_pf_num==0 && local_vf_num ==674 && local_vf_active==1) `toggle_tready(674)   
              else if (local_pf_num==0 && local_vf_num ==675 && local_vf_active==1) `toggle_tready(675)   
              else if (local_pf_num==0 && local_vf_num ==676 && local_vf_active==1) `toggle_tready(676)   
              else if (local_pf_num==0 && local_vf_num ==677 && local_vf_active==1) `toggle_tready(677)   
              else if (local_pf_num==0 && local_vf_num ==678 && local_vf_active==1) `toggle_tready(678)   
              else if (local_pf_num==0 && local_vf_num ==679 && local_vf_active==1) `toggle_tready(679)   
              else if (local_pf_num==0 && local_vf_num ==680 && local_vf_active==1) `toggle_tready(680)   
              else if (local_pf_num==0 && local_vf_num ==681 && local_vf_active==1) `toggle_tready(681)   
              else if (local_pf_num==0 && local_vf_num ==682 && local_vf_active==1) `toggle_tready(682)   
              else if (local_pf_num==0 && local_vf_num ==683 && local_vf_active==1) `toggle_tready(683)   
              else if (local_pf_num==0 && local_vf_num ==684 && local_vf_active==1) `toggle_tready(684)   
              else if (local_pf_num==0 && local_vf_num ==685 && local_vf_active==1) `toggle_tready(685)   
              else if (local_pf_num==0 && local_vf_num ==686 && local_vf_active==1) `toggle_tready(686)   
              else if (local_pf_num==0 && local_vf_num ==687 && local_vf_active==1) `toggle_tready(687)   
              else if (local_pf_num==0 && local_vf_num ==688 && local_vf_active==1) `toggle_tready(688)   
              else if (local_pf_num==0 && local_vf_num ==689 && local_vf_active==1) `toggle_tready(689)   
              else if (local_pf_num==0 && local_vf_num ==690 && local_vf_active==1) `toggle_tready(690)   
              else if (local_pf_num==0 && local_vf_num ==691 && local_vf_active==1) `toggle_tready(691)   
              else if (local_pf_num==0 && local_vf_num ==692 && local_vf_active==1) `toggle_tready(692)   
              else if (local_pf_num==0 && local_vf_num ==693 && local_vf_active==1) `toggle_tready(693)   
              else if (local_pf_num==0 && local_vf_num ==694 && local_vf_active==1) `toggle_tready(694)   
              else if (local_pf_num==0 && local_vf_num ==695 && local_vf_active==1) `toggle_tready(695)   
              else if (local_pf_num==0 && local_vf_num ==696 && local_vf_active==1) `toggle_tready(696)   
              else if (local_pf_num==0 && local_vf_num ==697 && local_vf_active==1) `toggle_tready(697)   
              else if (local_pf_num==0 && local_vf_num ==698 && local_vf_active==1) `toggle_tready(698)   
              else if (local_pf_num==0 && local_vf_num ==699 && local_vf_active==1) `toggle_tready(699)   
              else if (local_pf_num==0 && local_vf_num ==700 && local_vf_active==1) `toggle_tready(700)   
              else if (local_pf_num==0 && local_vf_num ==701 && local_vf_active==1) `toggle_tready(701)   
              else if (local_pf_num==0 && local_vf_num ==702 && local_vf_active==1) `toggle_tready(702)   
              else if (local_pf_num==0 && local_vf_num ==703 && local_vf_active==1) `toggle_tready(703)   
              else if (local_pf_num==0 && local_vf_num ==704 && local_vf_active==1) `toggle_tready(704)   
              else if (local_pf_num==0 && local_vf_num ==705 && local_vf_active==1) `toggle_tready(705)   
              else if (local_pf_num==0 && local_vf_num ==706 && local_vf_active==1) `toggle_tready(706)   
              else if (local_pf_num==0 && local_vf_num ==707 && local_vf_active==1) `toggle_tready(707)   
              else if (local_pf_num==0 && local_vf_num ==708 && local_vf_active==1) `toggle_tready(708)   
              else if (local_pf_num==0 && local_vf_num ==709 && local_vf_active==1) `toggle_tready(709)   
              else if (local_pf_num==0 && local_vf_num ==710 && local_vf_active==1) `toggle_tready(710)   
              else if (local_pf_num==0 && local_vf_num ==711 && local_vf_active==1) `toggle_tready(711)   
              else if (local_pf_num==0 && local_vf_num ==712 && local_vf_active==1) `toggle_tready(712)   
              else if (local_pf_num==0 && local_vf_num ==713 && local_vf_active==1) `toggle_tready(713)   
              else if (local_pf_num==0 && local_vf_num ==714 && local_vf_active==1) `toggle_tready(714)   
              else if (local_pf_num==0 && local_vf_num ==715 && local_vf_active==1) `toggle_tready(715)   
              else if (local_pf_num==0 && local_vf_num ==716 && local_vf_active==1) `toggle_tready(716)   
              else if (local_pf_num==0 && local_vf_num ==717 && local_vf_active==1) `toggle_tready(717)   
              else if (local_pf_num==0 && local_vf_num ==718 && local_vf_active==1) `toggle_tready(718)   
              else if (local_pf_num==0 && local_vf_num ==719 && local_vf_active==1) `toggle_tready(719)   
              else if (local_pf_num==0 && local_vf_num ==720 && local_vf_active==1) `toggle_tready(720)   
              else if (local_pf_num==0 && local_vf_num ==721 && local_vf_active==1) `toggle_tready(721)   
              else if (local_pf_num==0 && local_vf_num ==722 && local_vf_active==1) `toggle_tready(722)   
              else if (local_pf_num==0 && local_vf_num ==723 && local_vf_active==1) `toggle_tready(723)   
              else if (local_pf_num==0 && local_vf_num ==724 && local_vf_active==1) `toggle_tready(724)   
              else if (local_pf_num==0 && local_vf_num ==725 && local_vf_active==1) `toggle_tready(725)   
              else if (local_pf_num==0 && local_vf_num ==726 && local_vf_active==1) `toggle_tready(726)   
              else if (local_pf_num==0 && local_vf_num ==727 && local_vf_active==1) `toggle_tready(727)   
              else if (local_pf_num==0 && local_vf_num ==728 && local_vf_active==1) `toggle_tready(728)   
              else if (local_pf_num==0 && local_vf_num ==729 && local_vf_active==1) `toggle_tready(729)   
              else if (local_pf_num==0 && local_vf_num ==730 && local_vf_active==1) `toggle_tready(730)   
              else if (local_pf_num==0 && local_vf_num ==731 && local_vf_active==1) `toggle_tready(731)   
              else if (local_pf_num==0 && local_vf_num ==732 && local_vf_active==1) `toggle_tready(732)   
              else if (local_pf_num==0 && local_vf_num ==733 && local_vf_active==1) `toggle_tready(733)   
              else if (local_pf_num==0 && local_vf_num ==734 && local_vf_active==1) `toggle_tready(734)   
              else if (local_pf_num==0 && local_vf_num ==735 && local_vf_active==1) `toggle_tready(735)   
              else if (local_pf_num==0 && local_vf_num ==736 && local_vf_active==1) `toggle_tready(736)   
              else if (local_pf_num==0 && local_vf_num ==737 && local_vf_active==1) `toggle_tready(737)   
              else if (local_pf_num==0 && local_vf_num ==738 && local_vf_active==1) `toggle_tready(738)   
              else if (local_pf_num==0 && local_vf_num ==739 && local_vf_active==1) `toggle_tready(739)   
              else if (local_pf_num==0 && local_vf_num ==740 && local_vf_active==1) `toggle_tready(740)   
              else if (local_pf_num==0 && local_vf_num ==741 && local_vf_active==1) `toggle_tready(741)   
              else if (local_pf_num==0 && local_vf_num ==742 && local_vf_active==1) `toggle_tready(742)   
              else if (local_pf_num==0 && local_vf_num ==743 && local_vf_active==1) `toggle_tready(743)   
              else if (local_pf_num==0 && local_vf_num ==744 && local_vf_active==1) `toggle_tready(744)   
              else if (local_pf_num==0 && local_vf_num ==745 && local_vf_active==1) `toggle_tready(745)   
              else if (local_pf_num==0 && local_vf_num ==746 && local_vf_active==1) `toggle_tready(746)   
              else if (local_pf_num==0 && local_vf_num ==747 && local_vf_active==1) `toggle_tready(747)   
              else if (local_pf_num==0 && local_vf_num ==748 && local_vf_active==1) `toggle_tready(748)   
              else if (local_pf_num==0 && local_vf_num ==749 && local_vf_active==1) `toggle_tready(749)   
              else if (local_pf_num==0 && local_vf_num ==750 && local_vf_active==1) `toggle_tready(750)   
              else if (local_pf_num==0 && local_vf_num ==751 && local_vf_active==1) `toggle_tready(751)   
              else if (local_pf_num==0 && local_vf_num ==752 && local_vf_active==1) `toggle_tready(752)   
              else if (local_pf_num==0 && local_vf_num ==753 && local_vf_active==1) `toggle_tready(753)   
              else if (local_pf_num==0 && local_vf_num ==754 && local_vf_active==1) `toggle_tready(754)   
              else if (local_pf_num==0 && local_vf_num ==755 && local_vf_active==1) `toggle_tready(755)   
              else if (local_pf_num==0 && local_vf_num ==756 && local_vf_active==1) `toggle_tready(756)   
              else if (local_pf_num==0 && local_vf_num ==757 && local_vf_active==1) `toggle_tready(757)   
              else if (local_pf_num==0 && local_vf_num ==758 && local_vf_active==1) `toggle_tready(758)   
              else if (local_pf_num==0 && local_vf_num ==759 && local_vf_active==1) `toggle_tready(759)   
              else if (local_pf_num==0 && local_vf_num ==760 && local_vf_active==1) `toggle_tready(760)   
              else if (local_pf_num==0 && local_vf_num ==761 && local_vf_active==1) `toggle_tready(761)   
              else if (local_pf_num==0 && local_vf_num ==762 && local_vf_active==1) `toggle_tready(762)   
              else if (local_pf_num==0 && local_vf_num ==763 && local_vf_active==1) `toggle_tready(763)   
              else if (local_pf_num==0 && local_vf_num ==764 && local_vf_active==1) `toggle_tready(764)   
              else if (local_pf_num==0 && local_vf_num ==765 && local_vf_active==1) `toggle_tready(765)   
              else if (local_pf_num==0 && local_vf_num ==766 && local_vf_active==1) `toggle_tready(766)   
              else if (local_pf_num==0 && local_vf_num ==767 && local_vf_active==1) `toggle_tready(767)   
              else if (local_pf_num==0 && local_vf_num ==768 && local_vf_active==1) `toggle_tready(768)   
              else if (local_pf_num==0 && local_vf_num ==769 && local_vf_active==1) `toggle_tready(769)   
              else if (local_pf_num==0 && local_vf_num ==770 && local_vf_active==1) `toggle_tready(770)   
              else if (local_pf_num==0 && local_vf_num ==771 && local_vf_active==1) `toggle_tready(771)   
              else if (local_pf_num==0 && local_vf_num ==772 && local_vf_active==1) `toggle_tready(772)   
              else if (local_pf_num==0 && local_vf_num ==773 && local_vf_active==1) `toggle_tready(773)   
              else if (local_pf_num==0 && local_vf_num ==774 && local_vf_active==1) `toggle_tready(774)   
              else if (local_pf_num==0 && local_vf_num ==775 && local_vf_active==1) `toggle_tready(775)   
              else if (local_pf_num==0 && local_vf_num ==776 && local_vf_active==1) `toggle_tready(776)   
              else if (local_pf_num==0 && local_vf_num ==777 && local_vf_active==1) `toggle_tready(777)   
              else if (local_pf_num==0 && local_vf_num ==778 && local_vf_active==1) `toggle_tready(778)   
              else if (local_pf_num==0 && local_vf_num ==779 && local_vf_active==1) `toggle_tready(779)   
              else if (local_pf_num==0 && local_vf_num ==780 && local_vf_active==1) `toggle_tready(780)   
              else if (local_pf_num==0 && local_vf_num ==781 && local_vf_active==1) `toggle_tready(781)   
              else if (local_pf_num==0 && local_vf_num ==782 && local_vf_active==1) `toggle_tready(782)   
              else if (local_pf_num==0 && local_vf_num ==783 && local_vf_active==1) `toggle_tready(783)   
              else if (local_pf_num==0 && local_vf_num ==784 && local_vf_active==1) `toggle_tready(784)   
              else if (local_pf_num==0 && local_vf_num ==785 && local_vf_active==1) `toggle_tready(785)   
              else if (local_pf_num==0 && local_vf_num ==786 && local_vf_active==1) `toggle_tready(786)   
              else if (local_pf_num==0 && local_vf_num ==787 && local_vf_active==1) `toggle_tready(787)   
              else if (local_pf_num==0 && local_vf_num ==788 && local_vf_active==1) `toggle_tready(788)   
              else if (local_pf_num==0 && local_vf_num ==789 && local_vf_active==1) `toggle_tready(789)   
              else if (local_pf_num==0 && local_vf_num ==790 && local_vf_active==1) `toggle_tready(790)   
              else if (local_pf_num==0 && local_vf_num ==791 && local_vf_active==1) `toggle_tready(791)   
              else if (local_pf_num==0 && local_vf_num ==792 && local_vf_active==1) `toggle_tready(792)   
              else if (local_pf_num==0 && local_vf_num ==793 && local_vf_active==1) `toggle_tready(793)   
              else if (local_pf_num==0 && local_vf_num ==794 && local_vf_active==1) `toggle_tready(794)   
              else if (local_pf_num==0 && local_vf_num ==795 && local_vf_active==1) `toggle_tready(795)   
              else if (local_pf_num==0 && local_vf_num ==796 && local_vf_active==1) `toggle_tready(796)   
              else if (local_pf_num==0 && local_vf_num ==797 && local_vf_active==1) `toggle_tready(797)   
              else if (local_pf_num==0 && local_vf_num ==798 && local_vf_active==1) `toggle_tready(798)   
              else if (local_pf_num==0 && local_vf_num ==799 && local_vf_active==1) `toggle_tready(799)   
              else if (local_pf_num==0 && local_vf_num ==800 && local_vf_active==1) `toggle_tready(800)   
              else if (local_pf_num==0 && local_vf_num ==801 && local_vf_active==1) `toggle_tready(801)   
              else if (local_pf_num==0 && local_vf_num ==802 && local_vf_active==1) `toggle_tready(802)   
              else if (local_pf_num==0 && local_vf_num ==803 && local_vf_active==1) `toggle_tready(803)   
              else if (local_pf_num==0 && local_vf_num ==804 && local_vf_active==1) `toggle_tready(804)   
              else if (local_pf_num==0 && local_vf_num ==805 && local_vf_active==1) `toggle_tready(805)   
              else if (local_pf_num==0 && local_vf_num ==806 && local_vf_active==1) `toggle_tready(806)   
              else if (local_pf_num==0 && local_vf_num ==807 && local_vf_active==1) `toggle_tready(807)   
              else if (local_pf_num==0 && local_vf_num ==808 && local_vf_active==1) `toggle_tready(808)   
              else if (local_pf_num==0 && local_vf_num ==809 && local_vf_active==1) `toggle_tready(809)   
              else if (local_pf_num==0 && local_vf_num ==810 && local_vf_active==1) `toggle_tready(810)   
              else if (local_pf_num==0 && local_vf_num ==811 && local_vf_active==1) `toggle_tready(811)   
              else if (local_pf_num==0 && local_vf_num ==812 && local_vf_active==1) `toggle_tready(812)   
              else if (local_pf_num==0 && local_vf_num ==813 && local_vf_active==1) `toggle_tready(813)   
              else if (local_pf_num==0 && local_vf_num ==814 && local_vf_active==1) `toggle_tready(814)   
              else if (local_pf_num==0 && local_vf_num ==815 && local_vf_active==1) `toggle_tready(815)   
              else if (local_pf_num==0 && local_vf_num ==816 && local_vf_active==1) `toggle_tready(816)   
              else if (local_pf_num==0 && local_vf_num ==817 && local_vf_active==1) `toggle_tready(817)   
              else if (local_pf_num==0 && local_vf_num ==818 && local_vf_active==1) `toggle_tready(818)   
              else if (local_pf_num==0 && local_vf_num ==819 && local_vf_active==1) `toggle_tready(819)   
              else if (local_pf_num==0 && local_vf_num ==820 && local_vf_active==1) `toggle_tready(820)   
              else if (local_pf_num==0 && local_vf_num ==821 && local_vf_active==1) `toggle_tready(821)   
              else if (local_pf_num==0 && local_vf_num ==822 && local_vf_active==1) `toggle_tready(822)   
              else if (local_pf_num==0 && local_vf_num ==823 && local_vf_active==1) `toggle_tready(823)   
              else if (local_pf_num==0 && local_vf_num ==824 && local_vf_active==1) `toggle_tready(824)   
              else if (local_pf_num==0 && local_vf_num ==825 && local_vf_active==1) `toggle_tready(825)   
              else if (local_pf_num==0 && local_vf_num ==826 && local_vf_active==1) `toggle_tready(826)   
              else if (local_pf_num==0 && local_vf_num ==827 && local_vf_active==1) `toggle_tready(827)   
              else if (local_pf_num==0 && local_vf_num ==828 && local_vf_active==1) `toggle_tready(828)   
              else if (local_pf_num==0 && local_vf_num ==829 && local_vf_active==1) `toggle_tready(829)   
              else if (local_pf_num==0 && local_vf_num ==830 && local_vf_active==1) `toggle_tready(830)   
              else if (local_pf_num==0 && local_vf_num ==831 && local_vf_active==1) `toggle_tready(831)   
              else if (local_pf_num==0 && local_vf_num ==832 && local_vf_active==1) `toggle_tready(832)   
              else if (local_pf_num==0 && local_vf_num ==833 && local_vf_active==1) `toggle_tready(833)   
              else if (local_pf_num==0 && local_vf_num ==834 && local_vf_active==1) `toggle_tready(834)   
              else if (local_pf_num==0 && local_vf_num ==835 && local_vf_active==1) `toggle_tready(835)   
              else if (local_pf_num==0 && local_vf_num ==836 && local_vf_active==1) `toggle_tready(836)   
              else if (local_pf_num==0 && local_vf_num ==837 && local_vf_active==1) `toggle_tready(837)   
              else if (local_pf_num==0 && local_vf_num ==838 && local_vf_active==1) `toggle_tready(838)   
              else if (local_pf_num==0 && local_vf_num ==839 && local_vf_active==1) `toggle_tready(839)   
              else if (local_pf_num==0 && local_vf_num ==840 && local_vf_active==1) `toggle_tready(840)   
              else if (local_pf_num==0 && local_vf_num ==841 && local_vf_active==1) `toggle_tready(841)   
              else if (local_pf_num==0 && local_vf_num ==842 && local_vf_active==1) `toggle_tready(842)   
              else if (local_pf_num==0 && local_vf_num ==843 && local_vf_active==1) `toggle_tready(843)   
              else if (local_pf_num==0 && local_vf_num ==844 && local_vf_active==1) `toggle_tready(844)   
              else if (local_pf_num==0 && local_vf_num ==845 && local_vf_active==1) `toggle_tready(845)   
              else if (local_pf_num==0 && local_vf_num ==846 && local_vf_active==1) `toggle_tready(846)   
              else if (local_pf_num==0 && local_vf_num ==847 && local_vf_active==1) `toggle_tready(847)   
              else if (local_pf_num==0 && local_vf_num ==848 && local_vf_active==1) `toggle_tready(848)   
              else if (local_pf_num==0 && local_vf_num ==849 && local_vf_active==1) `toggle_tready(849)   
              else if (local_pf_num==0 && local_vf_num ==850 && local_vf_active==1) `toggle_tready(850)   
              else if (local_pf_num==0 && local_vf_num ==851 && local_vf_active==1) `toggle_tready(851)   
              else if (local_pf_num==0 && local_vf_num ==852 && local_vf_active==1) `toggle_tready(852)   
              else if (local_pf_num==0 && local_vf_num ==853 && local_vf_active==1) `toggle_tready(853)   
              else if (local_pf_num==0 && local_vf_num ==854 && local_vf_active==1) `toggle_tready(854)   
              else if (local_pf_num==0 && local_vf_num ==855 && local_vf_active==1) `toggle_tready(855)   
              else if (local_pf_num==0 && local_vf_num ==856 && local_vf_active==1) `toggle_tready(856)   
              else if (local_pf_num==0 && local_vf_num ==857 && local_vf_active==1) `toggle_tready(857)   
              else if (local_pf_num==0 && local_vf_num ==858 && local_vf_active==1) `toggle_tready(858)   
              else if (local_pf_num==0 && local_vf_num ==859 && local_vf_active==1) `toggle_tready(859)   
              else if (local_pf_num==0 && local_vf_num ==860 && local_vf_active==1) `toggle_tready(860)   
              else if (local_pf_num==0 && local_vf_num ==861 && local_vf_active==1) `toggle_tready(861)   
              else if (local_pf_num==0 && local_vf_num ==862 && local_vf_active==1) `toggle_tready(862)   
              else if (local_pf_num==0 && local_vf_num ==863 && local_vf_active==1) `toggle_tready(863)   
              else if (local_pf_num==0 && local_vf_num ==864 && local_vf_active==1) `toggle_tready(864)   
              else if (local_pf_num==0 && local_vf_num ==865 && local_vf_active==1) `toggle_tready(865)   
              else if (local_pf_num==0 && local_vf_num ==866 && local_vf_active==1) `toggle_tready(866)   
              else if (local_pf_num==0 && local_vf_num ==867 && local_vf_active==1) `toggle_tready(867)   
              else if (local_pf_num==0 && local_vf_num ==868 && local_vf_active==1) `toggle_tready(868)   
              else if (local_pf_num==0 && local_vf_num ==869 && local_vf_active==1) `toggle_tready(869)   
              else if (local_pf_num==0 && local_vf_num ==870 && local_vf_active==1) `toggle_tready(870)   
              else if (local_pf_num==0 && local_vf_num ==871 && local_vf_active==1) `toggle_tready(871)   
              else if (local_pf_num==0 && local_vf_num ==872 && local_vf_active==1) `toggle_tready(872)   
              else if (local_pf_num==0 && local_vf_num ==873 && local_vf_active==1) `toggle_tready(873)   
              else if (local_pf_num==0 && local_vf_num ==874 && local_vf_active==1) `toggle_tready(874)   
              else if (local_pf_num==0 && local_vf_num ==875 && local_vf_active==1) `toggle_tready(875)   
              else if (local_pf_num==0 && local_vf_num ==876 && local_vf_active==1) `toggle_tready(876)   
              else if (local_pf_num==0 && local_vf_num ==877 && local_vf_active==1) `toggle_tready(877)   
              else if (local_pf_num==0 && local_vf_num ==878 && local_vf_active==1) `toggle_tready(878)   
              else if (local_pf_num==0 && local_vf_num ==879 && local_vf_active==1) `toggle_tready(879)   
              else if (local_pf_num==0 && local_vf_num ==880 && local_vf_active==1) `toggle_tready(880)   
              else if (local_pf_num==0 && local_vf_num ==881 && local_vf_active==1) `toggle_tready(881)   
              else if (local_pf_num==0 && local_vf_num ==882 && local_vf_active==1) `toggle_tready(882)   
              else if (local_pf_num==0 && local_vf_num ==883 && local_vf_active==1) `toggle_tready(883)   
              else if (local_pf_num==0 && local_vf_num ==884 && local_vf_active==1) `toggle_tready(884)   
              else if (local_pf_num==0 && local_vf_num ==885 && local_vf_active==1) `toggle_tready(885)   
              else if (local_pf_num==0 && local_vf_num ==886 && local_vf_active==1) `toggle_tready(886)   
              else if (local_pf_num==0 && local_vf_num ==887 && local_vf_active==1) `toggle_tready(887)   
              else if (local_pf_num==0 && local_vf_num ==888 && local_vf_active==1) `toggle_tready(888)   
              else if (local_pf_num==0 && local_vf_num ==889 && local_vf_active==1) `toggle_tready(889)   
              else if (local_pf_num==0 && local_vf_num ==890 && local_vf_active==1) `toggle_tready(890)   
              else if (local_pf_num==0 && local_vf_num ==891 && local_vf_active==1) `toggle_tready(891)   
              else if (local_pf_num==0 && local_vf_num ==892 && local_vf_active==1) `toggle_tready(892)   
              else if (local_pf_num==0 && local_vf_num ==893 && local_vf_active==1) `toggle_tready(893)   
              else if (local_pf_num==0 && local_vf_num ==894 && local_vf_active==1) `toggle_tready(894)   
              else if (local_pf_num==0 && local_vf_num ==895 && local_vf_active==1) `toggle_tready(895)   
              else if (local_pf_num==0 && local_vf_num ==896 && local_vf_active==1) `toggle_tready(896)   
              else if (local_pf_num==0 && local_vf_num ==897 && local_vf_active==1) `toggle_tready(897)   
              else if (local_pf_num==0 && local_vf_num ==898 && local_vf_active==1) `toggle_tready(898)   
              else if (local_pf_num==0 && local_vf_num ==899 && local_vf_active==1) `toggle_tready(899)   
              else if (local_pf_num==0 && local_vf_num ==900 && local_vf_active==1) `toggle_tready(900)   
              else if (local_pf_num==0 && local_vf_num ==901 && local_vf_active==1) `toggle_tready(901)   
              else if (local_pf_num==0 && local_vf_num ==902 && local_vf_active==1) `toggle_tready(902)   
              else if (local_pf_num==0 && local_vf_num ==903 && local_vf_active==1) `toggle_tready(903)   
              else if (local_pf_num==0 && local_vf_num ==904 && local_vf_active==1) `toggle_tready(904)   
              else if (local_pf_num==0 && local_vf_num ==905 && local_vf_active==1) `toggle_tready(905)   
              else if (local_pf_num==0 && local_vf_num ==906 && local_vf_active==1) `toggle_tready(906)   
              else if (local_pf_num==0 && local_vf_num ==907 && local_vf_active==1) `toggle_tready(907)   
              else if (local_pf_num==0 && local_vf_num ==908 && local_vf_active==1) `toggle_tready(908)   
              else if (local_pf_num==0 && local_vf_num ==909 && local_vf_active==1) `toggle_tready(909)   
              else if (local_pf_num==0 && local_vf_num ==910 && local_vf_active==1) `toggle_tready(910)   
              else if (local_pf_num==0 && local_vf_num ==911 && local_vf_active==1) `toggle_tready(911)   
              else if (local_pf_num==0 && local_vf_num ==912 && local_vf_active==1) `toggle_tready(912)   
              else if (local_pf_num==0 && local_vf_num ==913 && local_vf_active==1) `toggle_tready(913)   
              else if (local_pf_num==0 && local_vf_num ==914 && local_vf_active==1) `toggle_tready(914)   
              else if (local_pf_num==0 && local_vf_num ==915 && local_vf_active==1) `toggle_tready(915)   
              else if (local_pf_num==0 && local_vf_num ==916 && local_vf_active==1) `toggle_tready(916)   
              else if (local_pf_num==0 && local_vf_num ==917 && local_vf_active==1) `toggle_tready(917)   
              else if (local_pf_num==0 && local_vf_num ==918 && local_vf_active==1) `toggle_tready(918)   
              else if (local_pf_num==0 && local_vf_num ==919 && local_vf_active==1) `toggle_tready(919)   
              else if (local_pf_num==0 && local_vf_num ==920 && local_vf_active==1) `toggle_tready(920)   
              else if (local_pf_num==0 && local_vf_num ==921 && local_vf_active==1) `toggle_tready(921)   
              else if (local_pf_num==0 && local_vf_num ==922 && local_vf_active==1) `toggle_tready(922)   
              else if (local_pf_num==0 && local_vf_num ==923 && local_vf_active==1) `toggle_tready(923)   
              else if (local_pf_num==0 && local_vf_num ==924 && local_vf_active==1) `toggle_tready(924)   
              else if (local_pf_num==0 && local_vf_num ==925 && local_vf_active==1) `toggle_tready(925)   
              else if (local_pf_num==0 && local_vf_num ==926 && local_vf_active==1) `toggle_tready(926)   
              else if (local_pf_num==0 && local_vf_num ==927 && local_vf_active==1) `toggle_tready(927)   
              else if (local_pf_num==0 && local_vf_num ==928 && local_vf_active==1) `toggle_tready(928)   
              else if (local_pf_num==0 && local_vf_num ==929 && local_vf_active==1) `toggle_tready(929)   
              else if (local_pf_num==0 && local_vf_num ==930 && local_vf_active==1) `toggle_tready(930)   
              else if (local_pf_num==0 && local_vf_num ==931 && local_vf_active==1) `toggle_tready(931)   
              else if (local_pf_num==0 && local_vf_num ==932 && local_vf_active==1) `toggle_tready(932)   
              else if (local_pf_num==0 && local_vf_num ==933 && local_vf_active==1) `toggle_tready(933)   
              else if (local_pf_num==0 && local_vf_num ==934 && local_vf_active==1) `toggle_tready(934)   
              else if (local_pf_num==0 && local_vf_num ==935 && local_vf_active==1) `toggle_tready(935)   
              else if (local_pf_num==0 && local_vf_num ==936 && local_vf_active==1) `toggle_tready(936)   
              else if (local_pf_num==0 && local_vf_num ==937 && local_vf_active==1) `toggle_tready(937)   
              else if (local_pf_num==0 && local_vf_num ==938 && local_vf_active==1) `toggle_tready(938)   
              else if (local_pf_num==0 && local_vf_num ==939 && local_vf_active==1) `toggle_tready(939)   
              else if (local_pf_num==0 && local_vf_num ==940 && local_vf_active==1) `toggle_tready(940)   
              else if (local_pf_num==0 && local_vf_num ==941 && local_vf_active==1) `toggle_tready(941)   
              else if (local_pf_num==0 && local_vf_num ==942 && local_vf_active==1) `toggle_tready(942)   
              else if (local_pf_num==0 && local_vf_num ==943 && local_vf_active==1) `toggle_tready(943)   
              else if (local_pf_num==0 && local_vf_num ==944 && local_vf_active==1) `toggle_tready(944)   
              else if (local_pf_num==0 && local_vf_num ==945 && local_vf_active==1) `toggle_tready(945)   
              else if (local_pf_num==0 && local_vf_num ==946 && local_vf_active==1) `toggle_tready(946)   
              else if (local_pf_num==0 && local_vf_num ==947 && local_vf_active==1) `toggle_tready(947)   
              else if (local_pf_num==0 && local_vf_num ==948 && local_vf_active==1) `toggle_tready(948)   
              else if (local_pf_num==0 && local_vf_num ==949 && local_vf_active==1) `toggle_tready(949)   
              else if (local_pf_num==0 && local_vf_num ==950 && local_vf_active==1) `toggle_tready(950)   
              else if (local_pf_num==0 && local_vf_num ==951 && local_vf_active==1) `toggle_tready(951)   
              else if (local_pf_num==0 && local_vf_num ==952 && local_vf_active==1) `toggle_tready(952)   
              else if (local_pf_num==0 && local_vf_num ==953 && local_vf_active==1) `toggle_tready(953)   
              else if (local_pf_num==0 && local_vf_num ==954 && local_vf_active==1) `toggle_tready(954)   
              else if (local_pf_num==0 && local_vf_num ==955 && local_vf_active==1) `toggle_tready(955)   
              else if (local_pf_num==0 && local_vf_num ==956 && local_vf_active==1) `toggle_tready(956)   
              else if (local_pf_num==0 && local_vf_num ==957 && local_vf_active==1) `toggle_tready(957)   
              else if (local_pf_num==0 && local_vf_num ==958 && local_vf_active==1) `toggle_tready(958)   
              else if (local_pf_num==0 && local_vf_num ==959 && local_vf_active==1) `toggle_tready(959)   
              else if (local_pf_num==0 && local_vf_num ==960 && local_vf_active==1) `toggle_tready(960)   
              else if (local_pf_num==0 && local_vf_num ==961 && local_vf_active==1) `toggle_tready(961)   
              else if (local_pf_num==0 && local_vf_num ==962 && local_vf_active==1) `toggle_tready(962)   
              else if (local_pf_num==0 && local_vf_num ==963 && local_vf_active==1) `toggle_tready(963)   
              else if (local_pf_num==0 && local_vf_num ==964 && local_vf_active==1) `toggle_tready(964)   
              else if (local_pf_num==0 && local_vf_num ==965 && local_vf_active==1) `toggle_tready(965)   
              else if (local_pf_num==0 && local_vf_num ==966 && local_vf_active==1) `toggle_tready(966)   
              else if (local_pf_num==0 && local_vf_num ==967 && local_vf_active==1) `toggle_tready(967)   
              else if (local_pf_num==0 && local_vf_num ==968 && local_vf_active==1) `toggle_tready(968)   
              else if (local_pf_num==0 && local_vf_num ==969 && local_vf_active==1) `toggle_tready(969)   
              else if (local_pf_num==0 && local_vf_num ==970 && local_vf_active==1) `toggle_tready(970)   
              else if (local_pf_num==0 && local_vf_num ==971 && local_vf_active==1) `toggle_tready(971)   
              else if (local_pf_num==0 && local_vf_num ==972 && local_vf_active==1) `toggle_tready(972)   
              else if (local_pf_num==0 && local_vf_num ==973 && local_vf_active==1) `toggle_tready(973)   
              else if (local_pf_num==0 && local_vf_num ==974 && local_vf_active==1) `toggle_tready(974)   
              else if (local_pf_num==0 && local_vf_num ==975 && local_vf_active==1) `toggle_tready(975)   
              else if (local_pf_num==0 && local_vf_num ==976 && local_vf_active==1) `toggle_tready(976)   
              else if (local_pf_num==0 && local_vf_num ==977 && local_vf_active==1) `toggle_tready(977)   
              else if (local_pf_num==0 && local_vf_num ==978 && local_vf_active==1) `toggle_tready(978)   
              else if (local_pf_num==0 && local_vf_num ==979 && local_vf_active==1) `toggle_tready(979)   
              else if (local_pf_num==0 && local_vf_num ==980 && local_vf_active==1) `toggle_tready(980)   
              else if (local_pf_num==0 && local_vf_num ==981 && local_vf_active==1) `toggle_tready(981)   
              else if (local_pf_num==0 && local_vf_num ==982 && local_vf_active==1) `toggle_tready(982)   
              else if (local_pf_num==0 && local_vf_num ==983 && local_vf_active==1) `toggle_tready(983)   
              else if (local_pf_num==0 && local_vf_num ==984 && local_vf_active==1) `toggle_tready(984)   
              else if (local_pf_num==0 && local_vf_num ==985 && local_vf_active==1) `toggle_tready(985)   
              else if (local_pf_num==0 && local_vf_num ==986 && local_vf_active==1) `toggle_tready(986)   
              else if (local_pf_num==0 && local_vf_num ==987 && local_vf_active==1) `toggle_tready(987)   
              else if (local_pf_num==0 && local_vf_num ==988 && local_vf_active==1) `toggle_tready(988)   
              else if (local_pf_num==0 && local_vf_num ==989 && local_vf_active==1) `toggle_tready(989)   
              else if (local_pf_num==0 && local_vf_num ==990 && local_vf_active==1) `toggle_tready(990)   
              else if (local_pf_num==0 && local_vf_num ==991 && local_vf_active==1) `toggle_tready(991)   
              else if (local_pf_num==0 && local_vf_num ==992 && local_vf_active==1) `toggle_tready(992)   
              else if (local_pf_num==0 && local_vf_num ==993 && local_vf_active==1) `toggle_tready(993)   
              else if (local_pf_num==0 && local_vf_num ==994 && local_vf_active==1) `toggle_tready(994)   
              else if (local_pf_num==0 && local_vf_num ==995 && local_vf_active==1) `toggle_tready(995)   
              else if (local_pf_num==0 && local_vf_num ==996 && local_vf_active==1) `toggle_tready(996)   
              else if (local_pf_num==0 && local_vf_num ==997 && local_vf_active==1) `toggle_tready(997)   
              else if (local_pf_num==0 && local_vf_num ==998 && local_vf_active==1) `toggle_tready(998)   
              else if (local_pf_num==0 && local_vf_num ==999 && local_vf_active==1) `toggle_tready(999)   
              else if (local_pf_num==0 && local_vf_num ==1000 && local_vf_active==1) `toggle_tready(1000)   
              else if (local_pf_num==0 && local_vf_num ==1001 && local_vf_active==1) `toggle_tready(1001)   
              else if (local_pf_num==0 && local_vf_num ==1002 && local_vf_active==1) `toggle_tready(1002)   
              else if (local_pf_num==0 && local_vf_num ==1003 && local_vf_active==1) `toggle_tready(1003)   
              else if (local_pf_num==0 && local_vf_num ==1004 && local_vf_active==1) `toggle_tready(1004)   
              else if (local_pf_num==0 && local_vf_num ==1005 && local_vf_active==1) `toggle_tready(1005)   
              else if (local_pf_num==0 && local_vf_num ==1006 && local_vf_active==1) `toggle_tready(1006)   
              else if (local_pf_num==0 && local_vf_num ==1007 && local_vf_active==1) `toggle_tready(1007)   
              else if (local_pf_num==0 && local_vf_num ==1008 && local_vf_active==1) `toggle_tready(1008)   
              else if (local_pf_num==0 && local_vf_num ==1009 && local_vf_active==1) `toggle_tready(1009)   
              else if (local_pf_num==0 && local_vf_num ==1010 && local_vf_active==1) `toggle_tready(1010)   
              else if (local_pf_num==0 && local_vf_num ==1011 && local_vf_active==1) `toggle_tready(1011)   
              else if (local_pf_num==0 && local_vf_num ==1012 && local_vf_active==1) `toggle_tready(1012)   
              else if (local_pf_num==0 && local_vf_num ==1013 && local_vf_active==1) `toggle_tready(1013)   
              else if (local_pf_num==0 && local_vf_num ==1014 && local_vf_active==1) `toggle_tready(1014)   
              else if (local_pf_num==0 && local_vf_num ==1015 && local_vf_active==1) `toggle_tready(1015)   
              else if (local_pf_num==0 && local_vf_num ==1016 && local_vf_active==1) `toggle_tready(1016)   
              else if (local_pf_num==0 && local_vf_num ==1017 && local_vf_active==1) `toggle_tready(1017)   
              else if (local_pf_num==0 && local_vf_num ==1018 && local_vf_active==1) `toggle_tready(1018)   
              else if (local_pf_num==0 && local_vf_num ==1019 && local_vf_active==1) `toggle_tready(1019)   
              else if (local_pf_num==0 && local_vf_num ==1020 && local_vf_active==1) `toggle_tready(1020)   
              else if (local_pf_num==0 && local_vf_num ==1021 && local_vf_active==1) `toggle_tready(1021)   
              else if (local_pf_num==0 && local_vf_num ==1022 && local_vf_active==1) `toggle_tready(1022)   
              else if (local_pf_num==0 && local_vf_num ==1023 && local_vf_active==1) `toggle_tready(1023)   
              else if (local_pf_num==0 && local_vf_num ==1024 && local_vf_active==1) `toggle_tready(1024)   
              else if (local_pf_num==0 && local_vf_num ==1025 && local_vf_active==1) `toggle_tready(1025)   
              else if (local_pf_num==0 && local_vf_num ==1026 && local_vf_active==1) `toggle_tready(1026)   
              else if (local_pf_num==0 && local_vf_num ==1027 && local_vf_active==1) `toggle_tready(1027)   
              else if (local_pf_num==0 && local_vf_num ==1028 && local_vf_active==1) `toggle_tready(1028)   
              else if (local_pf_num==0 && local_vf_num ==1029 && local_vf_active==1) `toggle_tready(1029)   
              else if (local_pf_num==0 && local_vf_num ==1030 && local_vf_active==1) `toggle_tready(1030)   
              else if (local_pf_num==0 && local_vf_num ==1031 && local_vf_active==1) `toggle_tready(1031)   
              else if (local_pf_num==0 && local_vf_num ==1032 && local_vf_active==1) `toggle_tready(1032)   
              else if (local_pf_num==0 && local_vf_num ==1033 && local_vf_active==1) `toggle_tready(1033)   
              else if (local_pf_num==0 && local_vf_num ==1034 && local_vf_active==1) `toggle_tready(1034)   
              else if (local_pf_num==0 && local_vf_num ==1035 && local_vf_active==1) `toggle_tready(1035)   
              else if (local_pf_num==0 && local_vf_num ==1036 && local_vf_active==1) `toggle_tready(1036)   
              else if (local_pf_num==0 && local_vf_num ==1037 && local_vf_active==1) `toggle_tready(1037)   
              else if (local_pf_num==0 && local_vf_num ==1038 && local_vf_active==1) `toggle_tready(1038)   
              else if (local_pf_num==0 && local_vf_num ==1039 && local_vf_active==1) `toggle_tready(1039)   
              else if (local_pf_num==0 && local_vf_num ==1040 && local_vf_active==1) `toggle_tready(1040)   
              else if (local_pf_num==0 && local_vf_num ==1041 && local_vf_active==1) `toggle_tready(1041)   
              else if (local_pf_num==0 && local_vf_num ==1042 && local_vf_active==1) `toggle_tready(1042)   
              else if (local_pf_num==0 && local_vf_num ==1043 && local_vf_active==1) `toggle_tready(1043)   
              else if (local_pf_num==0 && local_vf_num ==1044 && local_vf_active==1) `toggle_tready(1044)   
              else if (local_pf_num==0 && local_vf_num ==1045 && local_vf_active==1) `toggle_tready(1045)   
              else if (local_pf_num==0 && local_vf_num ==1046 && local_vf_active==1) `toggle_tready(1046)   
              else if (local_pf_num==0 && local_vf_num ==1047 && local_vf_active==1) `toggle_tready(1047)   
              else if (local_pf_num==0 && local_vf_num ==1048 && local_vf_active==1) `toggle_tready(1048)   
              else if (local_pf_num==0 && local_vf_num ==1049 && local_vf_active==1) `toggle_tready(1049)   
              else if (local_pf_num==0 && local_vf_num ==1050 && local_vf_active==1) `toggle_tready(1050)   
              else if (local_pf_num==0 && local_vf_num ==1051 && local_vf_active==1) `toggle_tready(1051)   
              else if (local_pf_num==0 && local_vf_num ==1052 && local_vf_active==1) `toggle_tready(1052)   
              else if (local_pf_num==0 && local_vf_num ==1053 && local_vf_active==1) `toggle_tready(1053)   
              else if (local_pf_num==0 && local_vf_num ==1054 && local_vf_active==1) `toggle_tready(1054)   
              else if (local_pf_num==0 && local_vf_num ==1055 && local_vf_active==1) `toggle_tready(1055)   
              else if (local_pf_num==0 && local_vf_num ==1056 && local_vf_active==1) `toggle_tready(1056)   
              else if (local_pf_num==0 && local_vf_num ==1057 && local_vf_active==1) `toggle_tready(1057)   
              else if (local_pf_num==0 && local_vf_num ==1058 && local_vf_active==1) `toggle_tready(1058)   
              else if (local_pf_num==0 && local_vf_num ==1059 && local_vf_active==1) `toggle_tready(1059)   
              else if (local_pf_num==0 && local_vf_num ==1060 && local_vf_active==1) `toggle_tready(1060)   
              else if (local_pf_num==0 && local_vf_num ==1061 && local_vf_active==1) `toggle_tready(1061)   
              else if (local_pf_num==0 && local_vf_num ==1062 && local_vf_active==1) `toggle_tready(1062)   
              else if (local_pf_num==0 && local_vf_num ==1063 && local_vf_active==1) `toggle_tready(1063)   
              else if (local_pf_num==0 && local_vf_num ==1064 && local_vf_active==1) `toggle_tready(1064)   
              else if (local_pf_num==0 && local_vf_num ==1065 && local_vf_active==1) `toggle_tready(1065)   
              else if (local_pf_num==0 && local_vf_num ==1066 && local_vf_active==1) `toggle_tready(1066)   
              else if (local_pf_num==0 && local_vf_num ==1067 && local_vf_active==1) `toggle_tready(1067)   
              else if (local_pf_num==0 && local_vf_num ==1068 && local_vf_active==1) `toggle_tready(1068)   
              else if (local_pf_num==0 && local_vf_num ==1069 && local_vf_active==1) `toggle_tready(1069)   
              else if (local_pf_num==0 && local_vf_num ==1070 && local_vf_active==1) `toggle_tready(1070)   
              else if (local_pf_num==0 && local_vf_num ==1071 && local_vf_active==1) `toggle_tready(1071)   
              else if (local_pf_num==0 && local_vf_num ==1072 && local_vf_active==1) `toggle_tready(1072)   
              else if (local_pf_num==0 && local_vf_num ==1073 && local_vf_active==1) `toggle_tready(1073)   
              else if (local_pf_num==0 && local_vf_num ==1074 && local_vf_active==1) `toggle_tready(1074)   
              else if (local_pf_num==0 && local_vf_num ==1075 && local_vf_active==1) `toggle_tready(1075)   
              else if (local_pf_num==0 && local_vf_num ==1076 && local_vf_active==1) `toggle_tready(1076)   
              else if (local_pf_num==0 && local_vf_num ==1077 && local_vf_active==1) `toggle_tready(1077)   
              else if (local_pf_num==0 && local_vf_num ==1078 && local_vf_active==1) `toggle_tready(1078)   
              else if (local_pf_num==0 && local_vf_num ==1079 && local_vf_active==1) `toggle_tready(1079)   
              else if (local_pf_num==0 && local_vf_num ==1080 && local_vf_active==1) `toggle_tready(1080)   
              else if (local_pf_num==0 && local_vf_num ==1081 && local_vf_active==1) `toggle_tready(1081)   
              else if (local_pf_num==0 && local_vf_num ==1082 && local_vf_active==1) `toggle_tready(1082)   
              else if (local_pf_num==0 && local_vf_num ==1083 && local_vf_active==1) `toggle_tready(1083)   
              else if (local_pf_num==0 && local_vf_num ==1084 && local_vf_active==1) `toggle_tready(1084)   
              else if (local_pf_num==0 && local_vf_num ==1085 && local_vf_active==1) `toggle_tready(1085)   
              else if (local_pf_num==0 && local_vf_num ==1086 && local_vf_active==1) `toggle_tready(1086)   
              else if (local_pf_num==0 && local_vf_num ==1087 && local_vf_active==1) `toggle_tready(1087)   
              else if (local_pf_num==0 && local_vf_num ==1088 && local_vf_active==1) `toggle_tready(1088)   
              else if (local_pf_num==0 && local_vf_num ==1089 && local_vf_active==1) `toggle_tready(1089)   
              else if (local_pf_num==0 && local_vf_num ==1090 && local_vf_active==1) `toggle_tready(1090)   
              else if (local_pf_num==0 && local_vf_num ==1091 && local_vf_active==1) `toggle_tready(1091)   
              else if (local_pf_num==0 && local_vf_num ==1092 && local_vf_active==1) `toggle_tready(1092)   
              else if (local_pf_num==0 && local_vf_num ==1093 && local_vf_active==1) `toggle_tready(1093)   
              else if (local_pf_num==0 && local_vf_num ==1094 && local_vf_active==1) `toggle_tready(1094)   
              else if (local_pf_num==0 && local_vf_num ==1095 && local_vf_active==1) `toggle_tready(1095)   
              else if (local_pf_num==0 && local_vf_num ==1096 && local_vf_active==1) `toggle_tready(1096)   
              else if (local_pf_num==0 && local_vf_num ==1097 && local_vf_active==1) `toggle_tready(1097)   
              else if (local_pf_num==0 && local_vf_num ==1098 && local_vf_active==1) `toggle_tready(1098)   
              else if (local_pf_num==0 && local_vf_num ==1099 && local_vf_active==1) `toggle_tready(1099)   
              else if (local_pf_num==0 && local_vf_num ==1100 && local_vf_active==1) `toggle_tready(1100)   
              else if (local_pf_num==0 && local_vf_num ==1101 && local_vf_active==1) `toggle_tready(1101)   
              else if (local_pf_num==0 && local_vf_num ==1102 && local_vf_active==1) `toggle_tready(1102)   
              else if (local_pf_num==0 && local_vf_num ==1103 && local_vf_active==1) `toggle_tready(1103)   
              else if (local_pf_num==0 && local_vf_num ==1104 && local_vf_active==1) `toggle_tready(1104)   
              else if (local_pf_num==0 && local_vf_num ==1105 && local_vf_active==1) `toggle_tready(1105)   
              else if (local_pf_num==0 && local_vf_num ==1106 && local_vf_active==1) `toggle_tready(1106)   
              else if (local_pf_num==0 && local_vf_num ==1107 && local_vf_active==1) `toggle_tready(1107)   
              else if (local_pf_num==0 && local_vf_num ==1108 && local_vf_active==1) `toggle_tready(1108)   
              else if (local_pf_num==0 && local_vf_num ==1109 && local_vf_active==1) `toggle_tready(1109)   
              else if (local_pf_num==0 && local_vf_num ==1110 && local_vf_active==1) `toggle_tready(1110)   
              else if (local_pf_num==0 && local_vf_num ==1111 && local_vf_active==1) `toggle_tready(1111)   
              else if (local_pf_num==0 && local_vf_num ==1112 && local_vf_active==1) `toggle_tready(1112)   
              else if (local_pf_num==0 && local_vf_num ==1113 && local_vf_active==1) `toggle_tready(1113)   
              else if (local_pf_num==0 && local_vf_num ==1114 && local_vf_active==1) `toggle_tready(1114)   
              else if (local_pf_num==0 && local_vf_num ==1115 && local_vf_active==1) `toggle_tready(1115)   
              else if (local_pf_num==0 && local_vf_num ==1116 && local_vf_active==1) `toggle_tready(1116)   
              else if (local_pf_num==0 && local_vf_num ==1117 && local_vf_active==1) `toggle_tready(1117)   
              else if (local_pf_num==0 && local_vf_num ==1118 && local_vf_active==1) `toggle_tready(1118)   
              else if (local_pf_num==0 && local_vf_num ==1119 && local_vf_active==1) `toggle_tready(1119)   
              else if (local_pf_num==0 && local_vf_num ==1120 && local_vf_active==1) `toggle_tready(1120)   
              else if (local_pf_num==0 && local_vf_num ==1121 && local_vf_active==1) `toggle_tready(1121)   
              else if (local_pf_num==0 && local_vf_num ==1122 && local_vf_active==1) `toggle_tready(1122)   
              else if (local_pf_num==0 && local_vf_num ==1123 && local_vf_active==1) `toggle_tready(1123)   
              else if (local_pf_num==0 && local_vf_num ==1124 && local_vf_active==1) `toggle_tready(1124)   
              else if (local_pf_num==0 && local_vf_num ==1125 && local_vf_active==1) `toggle_tready(1125)   
              else if (local_pf_num==0 && local_vf_num ==1126 && local_vf_active==1) `toggle_tready(1126)   
              else if (local_pf_num==0 && local_vf_num ==1127 && local_vf_active==1) `toggle_tready(1127)   
              else if (local_pf_num==0 && local_vf_num ==1128 && local_vf_active==1) `toggle_tready(1128)   
              else if (local_pf_num==0 && local_vf_num ==1129 && local_vf_active==1) `toggle_tready(1129)   
              else if (local_pf_num==0 && local_vf_num ==1130 && local_vf_active==1) `toggle_tready(1130)   
              else if (local_pf_num==0 && local_vf_num ==1131 && local_vf_active==1) `toggle_tready(1131)   
              else if (local_pf_num==0 && local_vf_num ==1132 && local_vf_active==1) `toggle_tready(1132)   
              else if (local_pf_num==0 && local_vf_num ==1133 && local_vf_active==1) `toggle_tready(1133)   
              else if (local_pf_num==0 && local_vf_num ==1134 && local_vf_active==1) `toggle_tready(1134)   
              else if (local_pf_num==0 && local_vf_num ==1135 && local_vf_active==1) `toggle_tready(1135)   
              else if (local_pf_num==0 && local_vf_num ==1136 && local_vf_active==1) `toggle_tready(1136)   
              else if (local_pf_num==0 && local_vf_num ==1137 && local_vf_active==1) `toggle_tready(1137)   
              else if (local_pf_num==0 && local_vf_num ==1138 && local_vf_active==1) `toggle_tready(1138)   
              else if (local_pf_num==0 && local_vf_num ==1139 && local_vf_active==1) `toggle_tready(1139)   
              else if (local_pf_num==0 && local_vf_num ==1140 && local_vf_active==1) `toggle_tready(1140)   
              else if (local_pf_num==0 && local_vf_num ==1141 && local_vf_active==1) `toggle_tready(1141)   
              else if (local_pf_num==0 && local_vf_num ==1142 && local_vf_active==1) `toggle_tready(1142)   
              else if (local_pf_num==0 && local_vf_num ==1143 && local_vf_active==1) `toggle_tready(1143)   
              else if (local_pf_num==0 && local_vf_num ==1144 && local_vf_active==1) `toggle_tready(1144)   
              else if (local_pf_num==0 && local_vf_num ==1145 && local_vf_active==1) `toggle_tready(1145)   
              else if (local_pf_num==0 && local_vf_num ==1146 && local_vf_active==1) `toggle_tready(1146)   
              else if (local_pf_num==0 && local_vf_num ==1147 && local_vf_active==1) `toggle_tready(1147)   
              else if (local_pf_num==0 && local_vf_num ==1148 && local_vf_active==1) `toggle_tready(1148)   
              else if (local_pf_num==0 && local_vf_num ==1149 && local_vf_active==1) `toggle_tready(1149)   
              else if (local_pf_num==0 && local_vf_num ==1150 && local_vf_active==1) `toggle_tready(1150)   
              else if (local_pf_num==0 && local_vf_num ==1151 && local_vf_active==1) `toggle_tready(1151)   
              else if (local_pf_num==0 && local_vf_num ==1152 && local_vf_active==1) `toggle_tready(1152)   
              else if (local_pf_num==0 && local_vf_num ==1153 && local_vf_active==1) `toggle_tready(1153)   
              else if (local_pf_num==0 && local_vf_num ==1154 && local_vf_active==1) `toggle_tready(1154)   
              else if (local_pf_num==0 && local_vf_num ==1155 && local_vf_active==1) `toggle_tready(1155)   
              else if (local_pf_num==0 && local_vf_num ==1156 && local_vf_active==1) `toggle_tready(1156)   
              else if (local_pf_num==0 && local_vf_num ==1157 && local_vf_active==1) `toggle_tready(1157)   
              else if (local_pf_num==0 && local_vf_num ==1158 && local_vf_active==1) `toggle_tready(1158)   
              else if (local_pf_num==0 && local_vf_num ==1159 && local_vf_active==1) `toggle_tready(1159)   
              else if (local_pf_num==0 && local_vf_num ==1160 && local_vf_active==1) `toggle_tready(1160)   
              else if (local_pf_num==0 && local_vf_num ==1161 && local_vf_active==1) `toggle_tready(1161)   
              else if (local_pf_num==0 && local_vf_num ==1162 && local_vf_active==1) `toggle_tready(1162)   
              else if (local_pf_num==0 && local_vf_num ==1163 && local_vf_active==1) `toggle_tready(1163)   
              else if (local_pf_num==0 && local_vf_num ==1164 && local_vf_active==1) `toggle_tready(1164)   
              else if (local_pf_num==0 && local_vf_num ==1165 && local_vf_active==1) `toggle_tready(1165)   
              else if (local_pf_num==0 && local_vf_num ==1166 && local_vf_active==1) `toggle_tready(1166)   
              else if (local_pf_num==0 && local_vf_num ==1167 && local_vf_active==1) `toggle_tready(1167)   
              else if (local_pf_num==0 && local_vf_num ==1168 && local_vf_active==1) `toggle_tready(1168)   
              else if (local_pf_num==0 && local_vf_num ==1169 && local_vf_active==1) `toggle_tready(1169)   
              else if (local_pf_num==0 && local_vf_num ==1170 && local_vf_active==1) `toggle_tready(1170)   
              else if (local_pf_num==0 && local_vf_num ==1171 && local_vf_active==1) `toggle_tready(1171)   
              else if (local_pf_num==0 && local_vf_num ==1172 && local_vf_active==1) `toggle_tready(1172)   
              else if (local_pf_num==0 && local_vf_num ==1173 && local_vf_active==1) `toggle_tready(1173)   
              else if (local_pf_num==0 && local_vf_num ==1174 && local_vf_active==1) `toggle_tready(1174)   
              else if (local_pf_num==0 && local_vf_num ==1175 && local_vf_active==1) `toggle_tready(1175)   
              else if (local_pf_num==0 && local_vf_num ==1176 && local_vf_active==1) `toggle_tready(1176)   
              else if (local_pf_num==0 && local_vf_num ==1177 && local_vf_active==1) `toggle_tready(1177)   
              else if (local_pf_num==0 && local_vf_num ==1178 && local_vf_active==1) `toggle_tready(1178)   
              else if (local_pf_num==0 && local_vf_num ==1179 && local_vf_active==1) `toggle_tready(1179)   
              else if (local_pf_num==0 && local_vf_num ==1180 && local_vf_active==1) `toggle_tready(1180)   
              else if (local_pf_num==0 && local_vf_num ==1181 && local_vf_active==1) `toggle_tready(1181)   
              else if (local_pf_num==0 && local_vf_num ==1182 && local_vf_active==1) `toggle_tready(1182)   
              else if (local_pf_num==0 && local_vf_num ==1183 && local_vf_active==1) `toggle_tready(1183)   
              else if (local_pf_num==0 && local_vf_num ==1184 && local_vf_active==1) `toggle_tready(1184)   
              else if (local_pf_num==0 && local_vf_num ==1185 && local_vf_active==1) `toggle_tready(1185)   
              else if (local_pf_num==0 && local_vf_num ==1186 && local_vf_active==1) `toggle_tready(1186)   
              else if (local_pf_num==0 && local_vf_num ==1187 && local_vf_active==1) `toggle_tready(1187)   
              else if (local_pf_num==0 && local_vf_num ==1188 && local_vf_active==1) `toggle_tready(1188)   
              else if (local_pf_num==0 && local_vf_num ==1189 && local_vf_active==1) `toggle_tready(1189)   
              else if (local_pf_num==0 && local_vf_num ==1190 && local_vf_active==1) `toggle_tready(1190)   
              else if (local_pf_num==0 && local_vf_num ==1191 && local_vf_active==1) `toggle_tready(1191)   
              else if (local_pf_num==0 && local_vf_num ==1192 && local_vf_active==1) `toggle_tready(1192)   
              else if (local_pf_num==0 && local_vf_num ==1193 && local_vf_active==1) `toggle_tready(1193)   
              else if (local_pf_num==0 && local_vf_num ==1194 && local_vf_active==1) `toggle_tready(1194)   
              else if (local_pf_num==0 && local_vf_num ==1195 && local_vf_active==1) `toggle_tready(1195)   
              else if (local_pf_num==0 && local_vf_num ==1196 && local_vf_active==1) `toggle_tready(1196)   
              else if (local_pf_num==0 && local_vf_num ==1197 && local_vf_active==1) `toggle_tready(1197)   
              else if (local_pf_num==0 && local_vf_num ==1198 && local_vf_active==1) `toggle_tready(1198)   
              else if (local_pf_num==0 && local_vf_num ==1199 && local_vf_active==1) `toggle_tready(1199)   
              else if (local_pf_num==0 && local_vf_num ==1200 && local_vf_active==1) `toggle_tready(1200)   
              else if (local_pf_num==0 && local_vf_num ==1201 && local_vf_active==1) `toggle_tready(1201)   
              else if (local_pf_num==0 && local_vf_num ==1202 && local_vf_active==1) `toggle_tready(1202)   
              else if (local_pf_num==0 && local_vf_num ==1203 && local_vf_active==1) `toggle_tready(1203)   
              else if (local_pf_num==0 && local_vf_num ==1204 && local_vf_active==1) `toggle_tready(1204)   
              else if (local_pf_num==0 && local_vf_num ==1205 && local_vf_active==1) `toggle_tready(1205)   
              else if (local_pf_num==0 && local_vf_num ==1206 && local_vf_active==1) `toggle_tready(1206)   
              else if (local_pf_num==0 && local_vf_num ==1207 && local_vf_active==1) `toggle_tready(1207)   
              else if (local_pf_num==0 && local_vf_num ==1208 && local_vf_active==1) `toggle_tready(1208)   
              else if (local_pf_num==0 && local_vf_num ==1209 && local_vf_active==1) `toggle_tready(1209)   
              else if (local_pf_num==0 && local_vf_num ==1210 && local_vf_active==1) `toggle_tready(1210)   
              else if (local_pf_num==0 && local_vf_num ==1211 && local_vf_active==1) `toggle_tready(1211)   
              else if (local_pf_num==0 && local_vf_num ==1212 && local_vf_active==1) `toggle_tready(1212)   
              else if (local_pf_num==0 && local_vf_num ==1213 && local_vf_active==1) `toggle_tready(1213)   
              else if (local_pf_num==0 && local_vf_num ==1214 && local_vf_active==1) `toggle_tready(1214)   
              else if (local_pf_num==0 && local_vf_num ==1215 && local_vf_active==1) `toggle_tready(1215)   
              else if (local_pf_num==0 && local_vf_num ==1216 && local_vf_active==1) `toggle_tready(1216)   
              else if (local_pf_num==0 && local_vf_num ==1217 && local_vf_active==1) `toggle_tready(1217)   
              else if (local_pf_num==0 && local_vf_num ==1218 && local_vf_active==1) `toggle_tready(1218)   
              else if (local_pf_num==0 && local_vf_num ==1219 && local_vf_active==1) `toggle_tready(1219)   
              else if (local_pf_num==0 && local_vf_num ==1220 && local_vf_active==1) `toggle_tready(1220)   
              else if (local_pf_num==0 && local_vf_num ==1221 && local_vf_active==1) `toggle_tready(1221)   
              else if (local_pf_num==0 && local_vf_num ==1222 && local_vf_active==1) `toggle_tready(1222)   
              else if (local_pf_num==0 && local_vf_num ==1223 && local_vf_active==1) `toggle_tready(1223)   
              else if (local_pf_num==0 && local_vf_num ==1224 && local_vf_active==1) `toggle_tready(1224)   
              else if (local_pf_num==0 && local_vf_num ==1225 && local_vf_active==1) `toggle_tready(1225)   
              else if (local_pf_num==0 && local_vf_num ==1226 && local_vf_active==1) `toggle_tready(1226)   
              else if (local_pf_num==0 && local_vf_num ==1227 && local_vf_active==1) `toggle_tready(1227)   
              else if (local_pf_num==0 && local_vf_num ==1228 && local_vf_active==1) `toggle_tready(1228)   
              else if (local_pf_num==0 && local_vf_num ==1229 && local_vf_active==1) `toggle_tready(1229)   
              else if (local_pf_num==0 && local_vf_num ==1230 && local_vf_active==1) `toggle_tready(1230)   
              else if (local_pf_num==0 && local_vf_num ==1231 && local_vf_active==1) `toggle_tready(1231)   
              else if (local_pf_num==0 && local_vf_num ==1232 && local_vf_active==1) `toggle_tready(1232)   
              else if (local_pf_num==0 && local_vf_num ==1233 && local_vf_active==1) `toggle_tready(1233)   
              else if (local_pf_num==0 && local_vf_num ==1234 && local_vf_active==1) `toggle_tready(1234)   
              else if (local_pf_num==0 && local_vf_num ==1235 && local_vf_active==1) `toggle_tready(1235)   
              else if (local_pf_num==0 && local_vf_num ==1236 && local_vf_active==1) `toggle_tready(1236)   
              else if (local_pf_num==0 && local_vf_num ==1237 && local_vf_active==1) `toggle_tready(1237)   
              else if (local_pf_num==0 && local_vf_num ==1238 && local_vf_active==1) `toggle_tready(1238)   
              else if (local_pf_num==0 && local_vf_num ==1239 && local_vf_active==1) `toggle_tready(1239)   
              else if (local_pf_num==0 && local_vf_num ==1240 && local_vf_active==1) `toggle_tready(1240)   
              else if (local_pf_num==0 && local_vf_num ==1241 && local_vf_active==1) `toggle_tready(1241)   
              else if (local_pf_num==0 && local_vf_num ==1242 && local_vf_active==1) `toggle_tready(1242)   
              else if (local_pf_num==0 && local_vf_num ==1243 && local_vf_active==1) `toggle_tready(1243)   
              else if (local_pf_num==0 && local_vf_num ==1244 && local_vf_active==1) `toggle_tready(1244)   
              else if (local_pf_num==0 && local_vf_num ==1245 && local_vf_active==1) `toggle_tready(1245)   
              else if (local_pf_num==0 && local_vf_num ==1246 && local_vf_active==1) `toggle_tready(1246)   
              else if (local_pf_num==0 && local_vf_num ==1247 && local_vf_active==1) `toggle_tready(1247)   
              else if (local_pf_num==0 && local_vf_num ==1248 && local_vf_active==1) `toggle_tready(1248)   
              else if (local_pf_num==0 && local_vf_num ==1249 && local_vf_active==1) `toggle_tready(1249)   
              else if (local_pf_num==0 && local_vf_num ==1250 && local_vf_active==1) `toggle_tready(1250)   
              else if (local_pf_num==0 && local_vf_num ==1251 && local_vf_active==1) `toggle_tready(1251)   
              else if (local_pf_num==0 && local_vf_num ==1252 && local_vf_active==1) `toggle_tready(1252)   
              else if (local_pf_num==0 && local_vf_num ==1253 && local_vf_active==1) `toggle_tready(1253)   
              else if (local_pf_num==0 && local_vf_num ==1254 && local_vf_active==1) `toggle_tready(1254)   
              else if (local_pf_num==0 && local_vf_num ==1255 && local_vf_active==1) `toggle_tready(1255)   
              else if (local_pf_num==0 && local_vf_num ==1256 && local_vf_active==1) `toggle_tready(1256)   
              else if (local_pf_num==0 && local_vf_num ==1257 && local_vf_active==1) `toggle_tready(1257)   
              else if (local_pf_num==0 && local_vf_num ==1258 && local_vf_active==1) `toggle_tready(1258)   
              else if (local_pf_num==0 && local_vf_num ==1259 && local_vf_active==1) `toggle_tready(1259)   
              else if (local_pf_num==0 && local_vf_num ==1260 && local_vf_active==1) `toggle_tready(1260)   
              else if (local_pf_num==0 && local_vf_num ==1261 && local_vf_active==1) `toggle_tready(1261)   
              else if (local_pf_num==0 && local_vf_num ==1262 && local_vf_active==1) `toggle_tready(1262)   
              else if (local_pf_num==0 && local_vf_num ==1263 && local_vf_active==1) `toggle_tready(1263)   
              else if (local_pf_num==0 && local_vf_num ==1264 && local_vf_active==1) `toggle_tready(1264)   
              else if (local_pf_num==0 && local_vf_num ==1265 && local_vf_active==1) `toggle_tready(1265)   
              else if (local_pf_num==0 && local_vf_num ==1266 && local_vf_active==1) `toggle_tready(1266)   
              else if (local_pf_num==0 && local_vf_num ==1267 && local_vf_active==1) `toggle_tready(1267)   
              else if (local_pf_num==0 && local_vf_num ==1268 && local_vf_active==1) `toggle_tready(1268)   
              else if (local_pf_num==0 && local_vf_num ==1269 && local_vf_active==1) `toggle_tready(1269)   
              else if (local_pf_num==0 && local_vf_num ==1270 && local_vf_active==1) `toggle_tready(1270)   
              else if (local_pf_num==0 && local_vf_num ==1271 && local_vf_active==1) `toggle_tready(1271)   
              else if (local_pf_num==0 && local_vf_num ==1272 && local_vf_active==1) `toggle_tready(1272)   
              else if (local_pf_num==0 && local_vf_num ==1273 && local_vf_active==1) `toggle_tready(1273)   
              else if (local_pf_num==0 && local_vf_num ==1274 && local_vf_active==1) `toggle_tready(1274)   
              else if (local_pf_num==0 && local_vf_num ==1275 && local_vf_active==1) `toggle_tready(1275)   
              else if (local_pf_num==0 && local_vf_num ==1276 && local_vf_active==1) `toggle_tready(1276)   
              else if (local_pf_num==0 && local_vf_num ==1277 && local_vf_active==1) `toggle_tready(1277)   
              else if (local_pf_num==0 && local_vf_num ==1278 && local_vf_active==1) `toggle_tready(1278)   
              else if (local_pf_num==0 && local_vf_num ==1279 && local_vf_active==1) `toggle_tready(1279)   
              else if (local_pf_num==0 && local_vf_num ==1280 && local_vf_active==1) `toggle_tready(1280)   
              else if (local_pf_num==0 && local_vf_num ==1281 && local_vf_active==1) `toggle_tready(1281)   
              else if (local_pf_num==0 && local_vf_num ==1282 && local_vf_active==1) `toggle_tready(1282)   
              else if (local_pf_num==0 && local_vf_num ==1283 && local_vf_active==1) `toggle_tready(1283)   
              else if (local_pf_num==0 && local_vf_num ==1284 && local_vf_active==1) `toggle_tready(1284)   
              else if (local_pf_num==0 && local_vf_num ==1285 && local_vf_active==1) `toggle_tready(1285)   
              else if (local_pf_num==0 && local_vf_num ==1286 && local_vf_active==1) `toggle_tready(1286)   
              else if (local_pf_num==0 && local_vf_num ==1287 && local_vf_active==1) `toggle_tready(1287)   
              else if (local_pf_num==0 && local_vf_num ==1288 && local_vf_active==1) `toggle_tready(1288)   
              else if (local_pf_num==0 && local_vf_num ==1289 && local_vf_active==1) `toggle_tready(1289)   
              else if (local_pf_num==0 && local_vf_num ==1290 && local_vf_active==1) `toggle_tready(1290)   
              else if (local_pf_num==0 && local_vf_num ==1291 && local_vf_active==1) `toggle_tready(1291)   
              else if (local_pf_num==0 && local_vf_num ==1292 && local_vf_active==1) `toggle_tready(1292)   
              else if (local_pf_num==0 && local_vf_num ==1293 && local_vf_active==1) `toggle_tready(1293)   
              else if (local_pf_num==0 && local_vf_num ==1294 && local_vf_active==1) `toggle_tready(1294)   
              else if (local_pf_num==0 && local_vf_num ==1295 && local_vf_active==1) `toggle_tready(1295)   
              else if (local_pf_num==0 && local_vf_num ==1296 && local_vf_active==1) `toggle_tready(1296)   
              else if (local_pf_num==0 && local_vf_num ==1297 && local_vf_active==1) `toggle_tready(1297)   
              else if (local_pf_num==0 && local_vf_num ==1298 && local_vf_active==1) `toggle_tready(1298)   
              else if (local_pf_num==0 && local_vf_num ==1299 && local_vf_active==1) `toggle_tready(1299)   
              else if (local_pf_num==0 && local_vf_num ==1300 && local_vf_active==1) `toggle_tready(1300)   
              else if (local_pf_num==0 && local_vf_num ==1301 && local_vf_active==1) `toggle_tready(1301)   
              else if (local_pf_num==0 && local_vf_num ==1302 && local_vf_active==1) `toggle_tready(1302)   
              else if (local_pf_num==0 && local_vf_num ==1303 && local_vf_active==1) `toggle_tready(1303)   
              else if (local_pf_num==0 && local_vf_num ==1304 && local_vf_active==1) `toggle_tready(1304)   
              else if (local_pf_num==0 && local_vf_num ==1305 && local_vf_active==1) `toggle_tready(1305)   
              else if (local_pf_num==0 && local_vf_num ==1306 && local_vf_active==1) `toggle_tready(1306)   
              else if (local_pf_num==0 && local_vf_num ==1307 && local_vf_active==1) `toggle_tready(1307)   
              else if (local_pf_num==0 && local_vf_num ==1308 && local_vf_active==1) `toggle_tready(1308)   
              else if (local_pf_num==0 && local_vf_num ==1309 && local_vf_active==1) `toggle_tready(1309)   
              else if (local_pf_num==0 && local_vf_num ==1310 && local_vf_active==1) `toggle_tready(1310)   
              else if (local_pf_num==0 && local_vf_num ==1311 && local_vf_active==1) `toggle_tready(1311)   
              else if (local_pf_num==0 && local_vf_num ==1312 && local_vf_active==1) `toggle_tready(1312)   
              else if (local_pf_num==0 && local_vf_num ==1313 && local_vf_active==1) `toggle_tready(1313)   
              else if (local_pf_num==0 && local_vf_num ==1314 && local_vf_active==1) `toggle_tready(1314)   
              else if (local_pf_num==0 && local_vf_num ==1315 && local_vf_active==1) `toggle_tready(1315)   
              else if (local_pf_num==0 && local_vf_num ==1316 && local_vf_active==1) `toggle_tready(1316)   
              else if (local_pf_num==0 && local_vf_num ==1317 && local_vf_active==1) `toggle_tready(1317)   
              else if (local_pf_num==0 && local_vf_num ==1318 && local_vf_active==1) `toggle_tready(1318)   
              else if (local_pf_num==0 && local_vf_num ==1319 && local_vf_active==1) `toggle_tready(1319)   
              else if (local_pf_num==0 && local_vf_num ==1320 && local_vf_active==1) `toggle_tready(1320)   
              else if (local_pf_num==0 && local_vf_num ==1321 && local_vf_active==1) `toggle_tready(1321)   
              else if (local_pf_num==0 && local_vf_num ==1322 && local_vf_active==1) `toggle_tready(1322)   
              else if (local_pf_num==0 && local_vf_num ==1323 && local_vf_active==1) `toggle_tready(1323)   
              else if (local_pf_num==0 && local_vf_num ==1324 && local_vf_active==1) `toggle_tready(1324)   
              else if (local_pf_num==0 && local_vf_num ==1325 && local_vf_active==1) `toggle_tready(1325)   
              else if (local_pf_num==0 && local_vf_num ==1326 && local_vf_active==1) `toggle_tready(1326)   
              else if (local_pf_num==0 && local_vf_num ==1327 && local_vf_active==1) `toggle_tready(1327)   
              else if (local_pf_num==0 && local_vf_num ==1328 && local_vf_active==1) `toggle_tready(1328)   
              else if (local_pf_num==0 && local_vf_num ==1329 && local_vf_active==1) `toggle_tready(1329)   
              else if (local_pf_num==0 && local_vf_num ==1330 && local_vf_active==1) `toggle_tready(1330)   
              else if (local_pf_num==0 && local_vf_num ==1331 && local_vf_active==1) `toggle_tready(1331)   
              else if (local_pf_num==0 && local_vf_num ==1332 && local_vf_active==1) `toggle_tready(1332)   
              else if (local_pf_num==0 && local_vf_num ==1333 && local_vf_active==1) `toggle_tready(1333)   
              else if (local_pf_num==0 && local_vf_num ==1334 && local_vf_active==1) `toggle_tready(1334)   
              else if (local_pf_num==0 && local_vf_num ==1335 && local_vf_active==1) `toggle_tready(1335)   
              else if (local_pf_num==0 && local_vf_num ==1336 && local_vf_active==1) `toggle_tready(1336)   
              else if (local_pf_num==0 && local_vf_num ==1337 && local_vf_active==1) `toggle_tready(1337)   
              else if (local_pf_num==0 && local_vf_num ==1338 && local_vf_active==1) `toggle_tready(1338)   
              else if (local_pf_num==0 && local_vf_num ==1339 && local_vf_active==1) `toggle_tready(1339)   
              else if (local_pf_num==0 && local_vf_num ==1340 && local_vf_active==1) `toggle_tready(1340)   
              else if (local_pf_num==0 && local_vf_num ==1341 && local_vf_active==1) `toggle_tready(1341)   
              else if (local_pf_num==0 && local_vf_num ==1342 && local_vf_active==1) `toggle_tready(1342)   
              else if (local_pf_num==0 && local_vf_num ==1343 && local_vf_active==1) `toggle_tready(1343)   
              else if (local_pf_num==0 && local_vf_num ==1344 && local_vf_active==1) `toggle_tready(1344)   
              else if (local_pf_num==0 && local_vf_num ==1345 && local_vf_active==1) `toggle_tready(1345)   
              else if (local_pf_num==0 && local_vf_num ==1346 && local_vf_active==1) `toggle_tready(1346)   
              else if (local_pf_num==0 && local_vf_num ==1347 && local_vf_active==1) `toggle_tready(1347)   
              else if (local_pf_num==0 && local_vf_num ==1348 && local_vf_active==1) `toggle_tready(1348)   
              else if (local_pf_num==0 && local_vf_num ==1349 && local_vf_active==1) `toggle_tready(1349)   
              else if (local_pf_num==0 && local_vf_num ==1350 && local_vf_active==1) `toggle_tready(1350)   
              else if (local_pf_num==0 && local_vf_num ==1351 && local_vf_active==1) `toggle_tready(1351)   
              else if (local_pf_num==0 && local_vf_num ==1352 && local_vf_active==1) `toggle_tready(1352)   
              else if (local_pf_num==0 && local_vf_num ==1353 && local_vf_active==1) `toggle_tready(1353)   
              else if (local_pf_num==0 && local_vf_num ==1354 && local_vf_active==1) `toggle_tready(1354)   
              else if (local_pf_num==0 && local_vf_num ==1355 && local_vf_active==1) `toggle_tready(1355)   
              else if (local_pf_num==0 && local_vf_num ==1356 && local_vf_active==1) `toggle_tready(1356)   
              else if (local_pf_num==0 && local_vf_num ==1357 && local_vf_active==1) `toggle_tready(1357)   
              else if (local_pf_num==0 && local_vf_num ==1358 && local_vf_active==1) `toggle_tready(1358)   
              else if (local_pf_num==0 && local_vf_num ==1359 && local_vf_active==1) `toggle_tready(1359)   
              else if (local_pf_num==0 && local_vf_num ==1360 && local_vf_active==1) `toggle_tready(1360)   
              else if (local_pf_num==0 && local_vf_num ==1361 && local_vf_active==1) `toggle_tready(1361)   
              else if (local_pf_num==0 && local_vf_num ==1362 && local_vf_active==1) `toggle_tready(1362)   
              else if (local_pf_num==0 && local_vf_num ==1363 && local_vf_active==1) `toggle_tready(1363)   
              else if (local_pf_num==0 && local_vf_num ==1364 && local_vf_active==1) `toggle_tready(1364)   
              else if (local_pf_num==0 && local_vf_num ==1365 && local_vf_active==1) `toggle_tready(1365)   
              else if (local_pf_num==0 && local_vf_num ==1366 && local_vf_active==1) `toggle_tready(1366)   
              else if (local_pf_num==0 && local_vf_num ==1367 && local_vf_active==1) `toggle_tready(1367)   
              else if (local_pf_num==0 && local_vf_num ==1368 && local_vf_active==1) `toggle_tready(1368)   
              else if (local_pf_num==0 && local_vf_num ==1369 && local_vf_active==1) `toggle_tready(1369)   
              else if (local_pf_num==0 && local_vf_num ==1370 && local_vf_active==1) `toggle_tready(1370)   
              else if (local_pf_num==0 && local_vf_num ==1371 && local_vf_active==1) `toggle_tready(1371)   
              else if (local_pf_num==0 && local_vf_num ==1372 && local_vf_active==1) `toggle_tready(1372)   
              else if (local_pf_num==0 && local_vf_num ==1373 && local_vf_active==1) `toggle_tready(1373)   
              else if (local_pf_num==0 && local_vf_num ==1374 && local_vf_active==1) `toggle_tready(1374)   
              else if (local_pf_num==0 && local_vf_num ==1375 && local_vf_active==1) `toggle_tready(1375)   
              else if (local_pf_num==0 && local_vf_num ==1376 && local_vf_active==1) `toggle_tready(1376)   
              else if (local_pf_num==0 && local_vf_num ==1377 && local_vf_active==1) `toggle_tready(1377)   
              else if (local_pf_num==0 && local_vf_num ==1378 && local_vf_active==1) `toggle_tready(1378)   
              else if (local_pf_num==0 && local_vf_num ==1379 && local_vf_active==1) `toggle_tready(1379)   
              else if (local_pf_num==0 && local_vf_num ==1380 && local_vf_active==1) `toggle_tready(1380)   
              else if (local_pf_num==0 && local_vf_num ==1381 && local_vf_active==1) `toggle_tready(1381)   
              else if (local_pf_num==0 && local_vf_num ==1382 && local_vf_active==1) `toggle_tready(1382)   
              else if (local_pf_num==0 && local_vf_num ==1383 && local_vf_active==1) `toggle_tready(1383)   
              else if (local_pf_num==0 && local_vf_num ==1384 && local_vf_active==1) `toggle_tready(1384)   
              else if (local_pf_num==0 && local_vf_num ==1385 && local_vf_active==1) `toggle_tready(1385)   
              else if (local_pf_num==0 && local_vf_num ==1386 && local_vf_active==1) `toggle_tready(1386)   
              else if (local_pf_num==0 && local_vf_num ==1387 && local_vf_active==1) `toggle_tready(1387)   
              else if (local_pf_num==0 && local_vf_num ==1388 && local_vf_active==1) `toggle_tready(1388)   
              else if (local_pf_num==0 && local_vf_num ==1389 && local_vf_active==1) `toggle_tready(1389)   
              else if (local_pf_num==0 && local_vf_num ==1390 && local_vf_active==1) `toggle_tready(1390)   
              else if (local_pf_num==0 && local_vf_num ==1391 && local_vf_active==1) `toggle_tready(1391)   
              else if (local_pf_num==0 && local_vf_num ==1392 && local_vf_active==1) `toggle_tready(1392)   
              else if (local_pf_num==0 && local_vf_num ==1393 && local_vf_active==1) `toggle_tready(1393)   
              else if (local_pf_num==0 && local_vf_num ==1394 && local_vf_active==1) `toggle_tready(1394)   
              else if (local_pf_num==0 && local_vf_num ==1395 && local_vf_active==1) `toggle_tready(1395)   
              else if (local_pf_num==0 && local_vf_num ==1396 && local_vf_active==1) `toggle_tready(1396)   
              else if (local_pf_num==0 && local_vf_num ==1397 && local_vf_active==1) `toggle_tready(1397)   
              else if (local_pf_num==0 && local_vf_num ==1398 && local_vf_active==1) `toggle_tready(1398)   
              else if (local_pf_num==0 && local_vf_num ==1399 && local_vf_active==1) `toggle_tready(1399)   
              else if (local_pf_num==0 && local_vf_num ==1400 && local_vf_active==1) `toggle_tready(1400)   
              else if (local_pf_num==0 && local_vf_num ==1401 && local_vf_active==1) `toggle_tready(1401)   
              else if (local_pf_num==0 && local_vf_num ==1402 && local_vf_active==1) `toggle_tready(1402)   
              else if (local_pf_num==0 && local_vf_num ==1403 && local_vf_active==1) `toggle_tready(1403)   
              else if (local_pf_num==0 && local_vf_num ==1404 && local_vf_active==1) `toggle_tready(1404)   
              else if (local_pf_num==0 && local_vf_num ==1405 && local_vf_active==1) `toggle_tready(1405)   
              else if (local_pf_num==0 && local_vf_num ==1406 && local_vf_active==1) `toggle_tready(1406)   
              else if (local_pf_num==0 && local_vf_num ==1407 && local_vf_active==1) `toggle_tready(1407)   
              else if (local_pf_num==0 && local_vf_num ==1408 && local_vf_active==1) `toggle_tready(1408)   
              else if (local_pf_num==0 && local_vf_num ==1409 && local_vf_active==1) `toggle_tready(1409)   
              else if (local_pf_num==0 && local_vf_num ==1410 && local_vf_active==1) `toggle_tready(1410)   
              else if (local_pf_num==0 && local_vf_num ==1411 && local_vf_active==1) `toggle_tready(1411)   
              else if (local_pf_num==0 && local_vf_num ==1412 && local_vf_active==1) `toggle_tready(1412)   
              else if (local_pf_num==0 && local_vf_num ==1413 && local_vf_active==1) `toggle_tready(1413)   
              else if (local_pf_num==0 && local_vf_num ==1414 && local_vf_active==1) `toggle_tready(1414)   
              else if (local_pf_num==0 && local_vf_num ==1415 && local_vf_active==1) `toggle_tready(1415)   
              else if (local_pf_num==0 && local_vf_num ==1416 && local_vf_active==1) `toggle_tready(1416)   
              else if (local_pf_num==0 && local_vf_num ==1417 && local_vf_active==1) `toggle_tready(1417)   
              else if (local_pf_num==0 && local_vf_num ==1418 && local_vf_active==1) `toggle_tready(1418)   
              else if (local_pf_num==0 && local_vf_num ==1419 && local_vf_active==1) `toggle_tready(1419)   
              else if (local_pf_num==0 && local_vf_num ==1420 && local_vf_active==1) `toggle_tready(1420)   
              else if (local_pf_num==0 && local_vf_num ==1421 && local_vf_active==1) `toggle_tready(1421)   
              else if (local_pf_num==0 && local_vf_num ==1422 && local_vf_active==1) `toggle_tready(1422)   
              else if (local_pf_num==0 && local_vf_num ==1423 && local_vf_active==1) `toggle_tready(1423)   
              else if (local_pf_num==0 && local_vf_num ==1424 && local_vf_active==1) `toggle_tready(1424)   
              else if (local_pf_num==0 && local_vf_num ==1425 && local_vf_active==1) `toggle_tready(1425)   
              else if (local_pf_num==0 && local_vf_num ==1426 && local_vf_active==1) `toggle_tready(1426)   
              else if (local_pf_num==0 && local_vf_num ==1427 && local_vf_active==1) `toggle_tready(1427)   
              else if (local_pf_num==0 && local_vf_num ==1428 && local_vf_active==1) `toggle_tready(1428)   
              else if (local_pf_num==0 && local_vf_num ==1429 && local_vf_active==1) `toggle_tready(1429)   
              else if (local_pf_num==0 && local_vf_num ==1430 && local_vf_active==1) `toggle_tready(1430)   
              else if (local_pf_num==0 && local_vf_num ==1431 && local_vf_active==1) `toggle_tready(1431)   
              else if (local_pf_num==0 && local_vf_num ==1432 && local_vf_active==1) `toggle_tready(1432)   
              else if (local_pf_num==0 && local_vf_num ==1433 && local_vf_active==1) `toggle_tready(1433)   
              else if (local_pf_num==0 && local_vf_num ==1434 && local_vf_active==1) `toggle_tready(1434)   
              else if (local_pf_num==0 && local_vf_num ==1435 && local_vf_active==1) `toggle_tready(1435)   
              else if (local_pf_num==0 && local_vf_num ==1436 && local_vf_active==1) `toggle_tready(1436)   
              else if (local_pf_num==0 && local_vf_num ==1437 && local_vf_active==1) `toggle_tready(1437)   
              else if (local_pf_num==0 && local_vf_num ==1438 && local_vf_active==1) `toggle_tready(1438)   
              else if (local_pf_num==0 && local_vf_num ==1439 && local_vf_active==1) `toggle_tready(1439)   
              else if (local_pf_num==0 && local_vf_num ==1440 && local_vf_active==1) `toggle_tready(1440)   
              else if (local_pf_num==0 && local_vf_num ==1441 && local_vf_active==1) `toggle_tready(1441)   
              else if (local_pf_num==0 && local_vf_num ==1442 && local_vf_active==1) `toggle_tready(1442)   
              else if (local_pf_num==0 && local_vf_num ==1443 && local_vf_active==1) `toggle_tready(1443)   
              else if (local_pf_num==0 && local_vf_num ==1444 && local_vf_active==1) `toggle_tready(1444)   
              else if (local_pf_num==0 && local_vf_num ==1445 && local_vf_active==1) `toggle_tready(1445)   
              else if (local_pf_num==0 && local_vf_num ==1446 && local_vf_active==1) `toggle_tready(1446)   
              else if (local_pf_num==0 && local_vf_num ==1447 && local_vf_active==1) `toggle_tready(1447)   
              else if (local_pf_num==0 && local_vf_num ==1448 && local_vf_active==1) `toggle_tready(1448)   
              else if (local_pf_num==0 && local_vf_num ==1449 && local_vf_active==1) `toggle_tready(1449)   
              else if (local_pf_num==0 && local_vf_num ==1450 && local_vf_active==1) `toggle_tready(1450)   
              else if (local_pf_num==0 && local_vf_num ==1451 && local_vf_active==1) `toggle_tready(1451)   
              else if (local_pf_num==0 && local_vf_num ==1452 && local_vf_active==1) `toggle_tready(1452)   
              else if (local_pf_num==0 && local_vf_num ==1453 && local_vf_active==1) `toggle_tready(1453)   
              else if (local_pf_num==0 && local_vf_num ==1454 && local_vf_active==1) `toggle_tready(1454)   
              else if (local_pf_num==0 && local_vf_num ==1455 && local_vf_active==1) `toggle_tready(1455)   
              else if (local_pf_num==0 && local_vf_num ==1456 && local_vf_active==1) `toggle_tready(1456)   
              else if (local_pf_num==0 && local_vf_num ==1457 && local_vf_active==1) `toggle_tready(1457)   
              else if (local_pf_num==0 && local_vf_num ==1458 && local_vf_active==1) `toggle_tready(1458)   
              else if (local_pf_num==0 && local_vf_num ==1459 && local_vf_active==1) `toggle_tready(1459)   
              else if (local_pf_num==0 && local_vf_num ==1460 && local_vf_active==1) `toggle_tready(1460)   
              else if (local_pf_num==0 && local_vf_num ==1461 && local_vf_active==1) `toggle_tready(1461)   
              else if (local_pf_num==0 && local_vf_num ==1462 && local_vf_active==1) `toggle_tready(1462)   
              else if (local_pf_num==0 && local_vf_num ==1463 && local_vf_active==1) `toggle_tready(1463)   
              else if (local_pf_num==0 && local_vf_num ==1464 && local_vf_active==1) `toggle_tready(1464)   
              else if (local_pf_num==0 && local_vf_num ==1465 && local_vf_active==1) `toggle_tready(1465)   
              else if (local_pf_num==0 && local_vf_num ==1466 && local_vf_active==1) `toggle_tready(1466)   
              else if (local_pf_num==0 && local_vf_num ==1467 && local_vf_active==1) `toggle_tready(1467)   
              else if (local_pf_num==0 && local_vf_num ==1468 && local_vf_active==1) `toggle_tready(1468)   
              else if (local_pf_num==0 && local_vf_num ==1469 && local_vf_active==1) `toggle_tready(1469)   
              else if (local_pf_num==0 && local_vf_num ==1470 && local_vf_active==1) `toggle_tready(1470)   
              else if (local_pf_num==0 && local_vf_num ==1471 && local_vf_active==1) `toggle_tready(1471)   
              else if (local_pf_num==0 && local_vf_num ==1472 && local_vf_active==1) `toggle_tready(1472)   
              else if (local_pf_num==0 && local_vf_num ==1473 && local_vf_active==1) `toggle_tready(1473)   
              else if (local_pf_num==0 && local_vf_num ==1474 && local_vf_active==1) `toggle_tready(1474)   
              else if (local_pf_num==0 && local_vf_num ==1475 && local_vf_active==1) `toggle_tready(1475)   
              else if (local_pf_num==0 && local_vf_num ==1476 && local_vf_active==1) `toggle_tready(1476)   
              else if (local_pf_num==0 && local_vf_num ==1477 && local_vf_active==1) `toggle_tready(1477)   
              else if (local_pf_num==0 && local_vf_num ==1478 && local_vf_active==1) `toggle_tready(1478)   
              else if (local_pf_num==0 && local_vf_num ==1479 && local_vf_active==1) `toggle_tready(1479)   
              else if (local_pf_num==0 && local_vf_num ==1480 && local_vf_active==1) `toggle_tready(1480)   
              else if (local_pf_num==0 && local_vf_num ==1481 && local_vf_active==1) `toggle_tready(1481)   
              else if (local_pf_num==0 && local_vf_num ==1482 && local_vf_active==1) `toggle_tready(1482)   
              else if (local_pf_num==0 && local_vf_num ==1483 && local_vf_active==1) `toggle_tready(1483)   
              else if (local_pf_num==0 && local_vf_num ==1484 && local_vf_active==1) `toggle_tready(1484)   
              else if (local_pf_num==0 && local_vf_num ==1485 && local_vf_active==1) `toggle_tready(1485)   
              else if (local_pf_num==0 && local_vf_num ==1486 && local_vf_active==1) `toggle_tready(1486)   
              else if (local_pf_num==0 && local_vf_num ==1487 && local_vf_active==1) `toggle_tready(1487)   
              else if (local_pf_num==0 && local_vf_num ==1488 && local_vf_active==1) `toggle_tready(1488)   
              else if (local_pf_num==0 && local_vf_num ==1489 && local_vf_active==1) `toggle_tready(1489)   
              else if (local_pf_num==0 && local_vf_num ==1490 && local_vf_active==1) `toggle_tready(1490)   
              else if (local_pf_num==0 && local_vf_num ==1491 && local_vf_active==1) `toggle_tready(1491)   
              else if (local_pf_num==0 && local_vf_num ==1492 && local_vf_active==1) `toggle_tready(1492)   
              else if (local_pf_num==0 && local_vf_num ==1493 && local_vf_active==1) `toggle_tready(1493)   
              else if (local_pf_num==0 && local_vf_num ==1494 && local_vf_active==1) `toggle_tready(1494)   
              else if (local_pf_num==0 && local_vf_num ==1495 && local_vf_active==1) `toggle_tready(1495)   
              else if (local_pf_num==0 && local_vf_num ==1496 && local_vf_active==1) `toggle_tready(1496)   
              else if (local_pf_num==0 && local_vf_num ==1497 && local_vf_active==1) `toggle_tready(1497)   
              else if (local_pf_num==0 && local_vf_num ==1498 && local_vf_active==1) `toggle_tready(1498)   
              else if (local_pf_num==0 && local_vf_num ==1499 && local_vf_active==1) `toggle_tready(1499)   
              else if (local_pf_num==0 && local_vf_num ==1500 && local_vf_active==1) `toggle_tready(1500)   
              else if (local_pf_num==0 && local_vf_num ==1501 && local_vf_active==1) `toggle_tready(1501)   
              else if (local_pf_num==0 && local_vf_num ==1502 && local_vf_active==1) `toggle_tready(1502)   
              else if (local_pf_num==0 && local_vf_num ==1503 && local_vf_active==1) `toggle_tready(1503)   
              else if (local_pf_num==0 && local_vf_num ==1504 && local_vf_active==1) `toggle_tready(1504)   
              else if (local_pf_num==0 && local_vf_num ==1505 && local_vf_active==1) `toggle_tready(1505)   
              else if (local_pf_num==0 && local_vf_num ==1506 && local_vf_active==1) `toggle_tready(1506)   
              else if (local_pf_num==0 && local_vf_num ==1507 && local_vf_active==1) `toggle_tready(1507)   
              else if (local_pf_num==0 && local_vf_num ==1508 && local_vf_active==1) `toggle_tready(1508)   
              else if (local_pf_num==0 && local_vf_num ==1509 && local_vf_active==1) `toggle_tready(1509)   
              else if (local_pf_num==0 && local_vf_num ==1510 && local_vf_active==1) `toggle_tready(1510)   
              else if (local_pf_num==0 && local_vf_num ==1511 && local_vf_active==1) `toggle_tready(1511)   
              else if (local_pf_num==0 && local_vf_num ==1512 && local_vf_active==1) `toggle_tready(1512)   
              else if (local_pf_num==0 && local_vf_num ==1513 && local_vf_active==1) `toggle_tready(1513)   
              else if (local_pf_num==0 && local_vf_num ==1514 && local_vf_active==1) `toggle_tready(1514)   
              else if (local_pf_num==0 && local_vf_num ==1515 && local_vf_active==1) `toggle_tready(1515)   
              else if (local_pf_num==0 && local_vf_num ==1516 && local_vf_active==1) `toggle_tready(1516)   
              else if (local_pf_num==0 && local_vf_num ==1517 && local_vf_active==1) `toggle_tready(1517)   
              else if (local_pf_num==0 && local_vf_num ==1518 && local_vf_active==1) `toggle_tready(1518)   
              else if (local_pf_num==0 && local_vf_num ==1519 && local_vf_active==1) `toggle_tready(1519)   
              else if (local_pf_num==0 && local_vf_num ==1520 && local_vf_active==1) `toggle_tready(1520)   
              else if (local_pf_num==0 && local_vf_num ==1521 && local_vf_active==1) `toggle_tready(1521)   
              else if (local_pf_num==0 && local_vf_num ==1522 && local_vf_active==1) `toggle_tready(1522)   
              else if (local_pf_num==0 && local_vf_num ==1523 && local_vf_active==1) `toggle_tready(1523)   
              else if (local_pf_num==0 && local_vf_num ==1524 && local_vf_active==1) `toggle_tready(1524)   
              else if (local_pf_num==0 && local_vf_num ==1525 && local_vf_active==1) `toggle_tready(1525)   
              else if (local_pf_num==0 && local_vf_num ==1526 && local_vf_active==1) `toggle_tready(1526)   
              else if (local_pf_num==0 && local_vf_num ==1527 && local_vf_active==1) `toggle_tready(1527)   
              else if (local_pf_num==0 && local_vf_num ==1528 && local_vf_active==1) `toggle_tready(1528)   
              else if (local_pf_num==0 && local_vf_num ==1529 && local_vf_active==1) `toggle_tready(1529)   
              else if (local_pf_num==0 && local_vf_num ==1530 && local_vf_active==1) `toggle_tready(1530)   
              else if (local_pf_num==0 && local_vf_num ==1531 && local_vf_active==1) `toggle_tready(1531)   
              else if (local_pf_num==0 && local_vf_num ==1532 && local_vf_active==1) `toggle_tready(1532)   
              else if (local_pf_num==0 && local_vf_num ==1533 && local_vf_active==1) `toggle_tready(1533)   
              else if (local_pf_num==0 && local_vf_num ==1534 && local_vf_active==1) `toggle_tready(1534)   
              else if (local_pf_num==0 && local_vf_num ==1535 && local_vf_active==1) `toggle_tready(1535)   
              else if (local_pf_num==0 && local_vf_num ==1536 && local_vf_active==1) `toggle_tready(1536)   
              else if (local_pf_num==0 && local_vf_num ==1537 && local_vf_active==1) `toggle_tready(1537)   
              else if (local_pf_num==0 && local_vf_num ==1538 && local_vf_active==1) `toggle_tready(1538)   
              else if (local_pf_num==0 && local_vf_num ==1539 && local_vf_active==1) `toggle_tready(1539)   
              else if (local_pf_num==0 && local_vf_num ==1540 && local_vf_active==1) `toggle_tready(1540)   
              else if (local_pf_num==0 && local_vf_num ==1541 && local_vf_active==1) `toggle_tready(1541)   
              else if (local_pf_num==0 && local_vf_num ==1542 && local_vf_active==1) `toggle_tready(1542)   
              else if (local_pf_num==0 && local_vf_num ==1543 && local_vf_active==1) `toggle_tready(1543)   
              else if (local_pf_num==0 && local_vf_num ==1544 && local_vf_active==1) `toggle_tready(1544)   
              else if (local_pf_num==0 && local_vf_num ==1545 && local_vf_active==1) `toggle_tready(1545)   
              else if (local_pf_num==0 && local_vf_num ==1546 && local_vf_active==1) `toggle_tready(1546)   
              else if (local_pf_num==0 && local_vf_num ==1547 && local_vf_active==1) `toggle_tready(1547)   
              else if (local_pf_num==0 && local_vf_num ==1548 && local_vf_active==1) `toggle_tready(1548)   
              else if (local_pf_num==0 && local_vf_num ==1549 && local_vf_active==1) `toggle_tready(1549)   
              else if (local_pf_num==0 && local_vf_num ==1550 && local_vf_active==1) `toggle_tready(1550)   
              else if (local_pf_num==0 && local_vf_num ==1551 && local_vf_active==1) `toggle_tready(1551)   
              else if (local_pf_num==0 && local_vf_num ==1552 && local_vf_active==1) `toggle_tready(1552)   
              else if (local_pf_num==0 && local_vf_num ==1553 && local_vf_active==1) `toggle_tready(1553)   
              else if (local_pf_num==0 && local_vf_num ==1554 && local_vf_active==1) `toggle_tready(1554)   
              else if (local_pf_num==0 && local_vf_num ==1555 && local_vf_active==1) `toggle_tready(1555)   
              else if (local_pf_num==0 && local_vf_num ==1556 && local_vf_active==1) `toggle_tready(1556)   
              else if (local_pf_num==0 && local_vf_num ==1557 && local_vf_active==1) `toggle_tready(1557)   
              else if (local_pf_num==0 && local_vf_num ==1558 && local_vf_active==1) `toggle_tready(1558)   
              else if (local_pf_num==0 && local_vf_num ==1559 && local_vf_active==1) `toggle_tready(1559)   
              else if (local_pf_num==0 && local_vf_num ==1560 && local_vf_active==1) `toggle_tready(1560)   
              else if (local_pf_num==0 && local_vf_num ==1561 && local_vf_active==1) `toggle_tready(1561)   
              else if (local_pf_num==0 && local_vf_num ==1562 && local_vf_active==1) `toggle_tready(1562)   
              else if (local_pf_num==0 && local_vf_num ==1563 && local_vf_active==1) `toggle_tready(1563)   
              else if (local_pf_num==0 && local_vf_num ==1564 && local_vf_active==1) `toggle_tready(1564)   
              else if (local_pf_num==0 && local_vf_num ==1565 && local_vf_active==1) `toggle_tready(1565)   
              else if (local_pf_num==0 && local_vf_num ==1566 && local_vf_active==1) `toggle_tready(1566)   
              else if (local_pf_num==0 && local_vf_num ==1567 && local_vf_active==1) `toggle_tready(1567)   
              else if (local_pf_num==0 && local_vf_num ==1568 && local_vf_active==1) `toggle_tready(1568)   
              else if (local_pf_num==0 && local_vf_num ==1569 && local_vf_active==1) `toggle_tready(1569)   
              else if (local_pf_num==0 && local_vf_num ==1570 && local_vf_active==1) `toggle_tready(1570)   
              else if (local_pf_num==0 && local_vf_num ==1571 && local_vf_active==1) `toggle_tready(1571)   
              else if (local_pf_num==0 && local_vf_num ==1572 && local_vf_active==1) `toggle_tready(1572)   
              else if (local_pf_num==0 && local_vf_num ==1573 && local_vf_active==1) `toggle_tready(1573)   
              else if (local_pf_num==0 && local_vf_num ==1574 && local_vf_active==1) `toggle_tready(1574)   
              else if (local_pf_num==0 && local_vf_num ==1575 && local_vf_active==1) `toggle_tready(1575)   
              else if (local_pf_num==0 && local_vf_num ==1576 && local_vf_active==1) `toggle_tready(1576)   
              else if (local_pf_num==0 && local_vf_num ==1577 && local_vf_active==1) `toggle_tready(1577)   
              else if (local_pf_num==0 && local_vf_num ==1578 && local_vf_active==1) `toggle_tready(1578)   
              else if (local_pf_num==0 && local_vf_num ==1579 && local_vf_active==1) `toggle_tready(1579)   
              else if (local_pf_num==0 && local_vf_num ==1580 && local_vf_active==1) `toggle_tready(1580)   
              else if (local_pf_num==0 && local_vf_num ==1581 && local_vf_active==1) `toggle_tready(1581)   
              else if (local_pf_num==0 && local_vf_num ==1582 && local_vf_active==1) `toggle_tready(1582)   
              else if (local_pf_num==0 && local_vf_num ==1583 && local_vf_active==1) `toggle_tready(1583)   
              else if (local_pf_num==0 && local_vf_num ==1584 && local_vf_active==1) `toggle_tready(1584)   
              else if (local_pf_num==0 && local_vf_num ==1585 && local_vf_active==1) `toggle_tready(1585)   
              else if (local_pf_num==0 && local_vf_num ==1586 && local_vf_active==1) `toggle_tready(1586)   
              else if (local_pf_num==0 && local_vf_num ==1587 && local_vf_active==1) `toggle_tready(1587)   
              else if (local_pf_num==0 && local_vf_num ==1588 && local_vf_active==1) `toggle_tready(1588)   
              else if (local_pf_num==0 && local_vf_num ==1589 && local_vf_active==1) `toggle_tready(1589)   
              else if (local_pf_num==0 && local_vf_num ==1590 && local_vf_active==1) `toggle_tready(1590)   
              else if (local_pf_num==0 && local_vf_num ==1591 && local_vf_active==1) `toggle_tready(1591)   
              else if (local_pf_num==0 && local_vf_num ==1592 && local_vf_active==1) `toggle_tready(1592)   
              else if (local_pf_num==0 && local_vf_num ==1593 && local_vf_active==1) `toggle_tready(1593)   
              else if (local_pf_num==0 && local_vf_num ==1594 && local_vf_active==1) `toggle_tready(1594)   
              else if (local_pf_num==0 && local_vf_num ==1595 && local_vf_active==1) `toggle_tready(1595)   
              else if (local_pf_num==0 && local_vf_num ==1596 && local_vf_active==1) `toggle_tready(1596)   
              else if (local_pf_num==0 && local_vf_num ==1597 && local_vf_active==1) `toggle_tready(1597)   
              else if (local_pf_num==0 && local_vf_num ==1598 && local_vf_active==1) `toggle_tready(1598)   
              else if (local_pf_num==0 && local_vf_num ==1599 && local_vf_active==1) `toggle_tready(1599)   
              else if (local_pf_num==0 && local_vf_num ==1600 && local_vf_active==1) `toggle_tready(1600)   
              else if (local_pf_num==0 && local_vf_num ==1601 && local_vf_active==1) `toggle_tready(1601)   
              else if (local_pf_num==0 && local_vf_num ==1602 && local_vf_active==1) `toggle_tready(1602)   
              else if (local_pf_num==0 && local_vf_num ==1603 && local_vf_active==1) `toggle_tready(1603)   
              else if (local_pf_num==0 && local_vf_num ==1604 && local_vf_active==1) `toggle_tready(1604)   
              else if (local_pf_num==0 && local_vf_num ==1605 && local_vf_active==1) `toggle_tready(1605)   
              else if (local_pf_num==0 && local_vf_num ==1606 && local_vf_active==1) `toggle_tready(1606)   
              else if (local_pf_num==0 && local_vf_num ==1607 && local_vf_active==1) `toggle_tready(1607)   
              else if (local_pf_num==0 && local_vf_num ==1608 && local_vf_active==1) `toggle_tready(1608)   
              else if (local_pf_num==0 && local_vf_num ==1609 && local_vf_active==1) `toggle_tready(1609)   
              else if (local_pf_num==0 && local_vf_num ==1610 && local_vf_active==1) `toggle_tready(1610)   
              else if (local_pf_num==0 && local_vf_num ==1611 && local_vf_active==1) `toggle_tready(1611)   
              else if (local_pf_num==0 && local_vf_num ==1612 && local_vf_active==1) `toggle_tready(1612)   
              else if (local_pf_num==0 && local_vf_num ==1613 && local_vf_active==1) `toggle_tready(1613)   
              else if (local_pf_num==0 && local_vf_num ==1614 && local_vf_active==1) `toggle_tready(1614)   
              else if (local_pf_num==0 && local_vf_num ==1615 && local_vf_active==1) `toggle_tready(1615)   
              else if (local_pf_num==0 && local_vf_num ==1616 && local_vf_active==1) `toggle_tready(1616)   
              else if (local_pf_num==0 && local_vf_num ==1617 && local_vf_active==1) `toggle_tready(1617)   
              else if (local_pf_num==0 && local_vf_num ==1618 && local_vf_active==1) `toggle_tready(1618)   
              else if (local_pf_num==0 && local_vf_num ==1619 && local_vf_active==1) `toggle_tready(1619)   
              else if (local_pf_num==0 && local_vf_num ==1620 && local_vf_active==1) `toggle_tready(1620)   
              else if (local_pf_num==0 && local_vf_num ==1621 && local_vf_active==1) `toggle_tready(1621)   
              else if (local_pf_num==0 && local_vf_num ==1622 && local_vf_active==1) `toggle_tready(1622)   
              else if (local_pf_num==0 && local_vf_num ==1623 && local_vf_active==1) `toggle_tready(1623)   
              else if (local_pf_num==0 && local_vf_num ==1624 && local_vf_active==1) `toggle_tready(1624)   
              else if (local_pf_num==0 && local_vf_num ==1625 && local_vf_active==1) `toggle_tready(1625)   
              else if (local_pf_num==0 && local_vf_num ==1626 && local_vf_active==1) `toggle_tready(1626)   
              else if (local_pf_num==0 && local_vf_num ==1627 && local_vf_active==1) `toggle_tready(1627)   
              else if (local_pf_num==0 && local_vf_num ==1628 && local_vf_active==1) `toggle_tready(1628)   
              else if (local_pf_num==0 && local_vf_num ==1629 && local_vf_active==1) `toggle_tready(1629)   
              else if (local_pf_num==0 && local_vf_num ==1630 && local_vf_active==1) `toggle_tready(1630)   
              else if (local_pf_num==0 && local_vf_num ==1631 && local_vf_active==1) `toggle_tready(1631)   
              else if (local_pf_num==0 && local_vf_num ==1632 && local_vf_active==1) `toggle_tready(1632)   
              else if (local_pf_num==0 && local_vf_num ==1633 && local_vf_active==1) `toggle_tready(1633)   
              else if (local_pf_num==0 && local_vf_num ==1634 && local_vf_active==1) `toggle_tready(1634)   
              else if (local_pf_num==0 && local_vf_num ==1635 && local_vf_active==1) `toggle_tready(1635)   
              else if (local_pf_num==0 && local_vf_num ==1636 && local_vf_active==1) `toggle_tready(1636)   
              else if (local_pf_num==0 && local_vf_num ==1637 && local_vf_active==1) `toggle_tready(1637)   
              else if (local_pf_num==0 && local_vf_num ==1638 && local_vf_active==1) `toggle_tready(1638)   
              else if (local_pf_num==0 && local_vf_num ==1639 && local_vf_active==1) `toggle_tready(1639)   
              else if (local_pf_num==0 && local_vf_num ==1640 && local_vf_active==1) `toggle_tready(1640)   
              else if (local_pf_num==0 && local_vf_num ==1641 && local_vf_active==1) `toggle_tready(1641)   
              else if (local_pf_num==0 && local_vf_num ==1642 && local_vf_active==1) `toggle_tready(1642)   
              else if (local_pf_num==0 && local_vf_num ==1643 && local_vf_active==1) `toggle_tready(1643)   
              else if (local_pf_num==0 && local_vf_num ==1644 && local_vf_active==1) `toggle_tready(1644)   
              else if (local_pf_num==0 && local_vf_num ==1645 && local_vf_active==1) `toggle_tready(1645)   
              else if (local_pf_num==0 && local_vf_num ==1646 && local_vf_active==1) `toggle_tready(1646)   
              else if (local_pf_num==0 && local_vf_num ==1647 && local_vf_active==1) `toggle_tready(1647)   
              else if (local_pf_num==0 && local_vf_num ==1648 && local_vf_active==1) `toggle_tready(1648)   
              else if (local_pf_num==0 && local_vf_num ==1649 && local_vf_active==1) `toggle_tready(1649)   
              else if (local_pf_num==0 && local_vf_num ==1650 && local_vf_active==1) `toggle_tready(1650)   
              else if (local_pf_num==0 && local_vf_num ==1651 && local_vf_active==1) `toggle_tready(1651)   
              else if (local_pf_num==0 && local_vf_num ==1652 && local_vf_active==1) `toggle_tready(1652)   
              else if (local_pf_num==0 && local_vf_num ==1653 && local_vf_active==1) `toggle_tready(1653)   
              else if (local_pf_num==0 && local_vf_num ==1654 && local_vf_active==1) `toggle_tready(1654)   
              else if (local_pf_num==0 && local_vf_num ==1655 && local_vf_active==1) `toggle_tready(1655)   
              else if (local_pf_num==0 && local_vf_num ==1656 && local_vf_active==1) `toggle_tready(1656)   
              else if (local_pf_num==0 && local_vf_num ==1657 && local_vf_active==1) `toggle_tready(1657)   
              else if (local_pf_num==0 && local_vf_num ==1658 && local_vf_active==1) `toggle_tready(1658)   
              else if (local_pf_num==0 && local_vf_num ==1659 && local_vf_active==1) `toggle_tready(1659)   
              else if (local_pf_num==0 && local_vf_num ==1660 && local_vf_active==1) `toggle_tready(1660)   
              else if (local_pf_num==0 && local_vf_num ==1661 && local_vf_active==1) `toggle_tready(1661)   
              else if (local_pf_num==0 && local_vf_num ==1662 && local_vf_active==1) `toggle_tready(1662)   
              else if (local_pf_num==0 && local_vf_num ==1663 && local_vf_active==1) `toggle_tready(1663)   
              else if (local_pf_num==0 && local_vf_num ==1664 && local_vf_active==1) `toggle_tready(1664)   
              else if (local_pf_num==0 && local_vf_num ==1665 && local_vf_active==1) `toggle_tready(1665)   
              else if (local_pf_num==0 && local_vf_num ==1666 && local_vf_active==1) `toggle_tready(1666)   
              else if (local_pf_num==0 && local_vf_num ==1667 && local_vf_active==1) `toggle_tready(1667)   
              else if (local_pf_num==0 && local_vf_num ==1668 && local_vf_active==1) `toggle_tready(1668)   
              else if (local_pf_num==0 && local_vf_num ==1669 && local_vf_active==1) `toggle_tready(1669)   
              else if (local_pf_num==0 && local_vf_num ==1670 && local_vf_active==1) `toggle_tready(1670)   
              else if (local_pf_num==0 && local_vf_num ==1671 && local_vf_active==1) `toggle_tready(1671)   
              else if (local_pf_num==0 && local_vf_num ==1672 && local_vf_active==1) `toggle_tready(1672)   
              else if (local_pf_num==0 && local_vf_num ==1673 && local_vf_active==1) `toggle_tready(1673)   
              else if (local_pf_num==0 && local_vf_num ==1674 && local_vf_active==1) `toggle_tready(1674)   
              else if (local_pf_num==0 && local_vf_num ==1675 && local_vf_active==1) `toggle_tready(1675)   
              else if (local_pf_num==0 && local_vf_num ==1676 && local_vf_active==1) `toggle_tready(1676)   
              else if (local_pf_num==0 && local_vf_num ==1677 && local_vf_active==1) `toggle_tready(1677)   
              else if (local_pf_num==0 && local_vf_num ==1678 && local_vf_active==1) `toggle_tready(1678)   
              else if (local_pf_num==0 && local_vf_num ==1679 && local_vf_active==1) `toggle_tready(1679)   
              else if (local_pf_num==0 && local_vf_num ==1680 && local_vf_active==1) `toggle_tready(1680)   
              else if (local_pf_num==0 && local_vf_num ==1681 && local_vf_active==1) `toggle_tready(1681)   
              else if (local_pf_num==0 && local_vf_num ==1682 && local_vf_active==1) `toggle_tready(1682)   
              else if (local_pf_num==0 && local_vf_num ==1683 && local_vf_active==1) `toggle_tready(1683)   
              else if (local_pf_num==0 && local_vf_num ==1684 && local_vf_active==1) `toggle_tready(1684)   
              else if (local_pf_num==0 && local_vf_num ==1685 && local_vf_active==1) `toggle_tready(1685)   
              else if (local_pf_num==0 && local_vf_num ==1686 && local_vf_active==1) `toggle_tready(1686)   
              else if (local_pf_num==0 && local_vf_num ==1687 && local_vf_active==1) `toggle_tready(1687)   
              else if (local_pf_num==0 && local_vf_num ==1688 && local_vf_active==1) `toggle_tready(1688)   
              else if (local_pf_num==0 && local_vf_num ==1689 && local_vf_active==1) `toggle_tready(1689)   
              else if (local_pf_num==0 && local_vf_num ==1690 && local_vf_active==1) `toggle_tready(1690)   
              else if (local_pf_num==0 && local_vf_num ==1691 && local_vf_active==1) `toggle_tready(1691)   
              else if (local_pf_num==0 && local_vf_num ==1692 && local_vf_active==1) `toggle_tready(1692)   
              else if (local_pf_num==0 && local_vf_num ==1693 && local_vf_active==1) `toggle_tready(1693)   
              else if (local_pf_num==0 && local_vf_num ==1694 && local_vf_active==1) `toggle_tready(1694)   
              else if (local_pf_num==0 && local_vf_num ==1695 && local_vf_active==1) `toggle_tready(1695)   
              else if (local_pf_num==0 && local_vf_num ==1696 && local_vf_active==1) `toggle_tready(1696)   
              else if (local_pf_num==0 && local_vf_num ==1697 && local_vf_active==1) `toggle_tready(1697)   
              else if (local_pf_num==0 && local_vf_num ==1698 && local_vf_active==1) `toggle_tready(1698)   
              else if (local_pf_num==0 && local_vf_num ==1699 && local_vf_active==1) `toggle_tready(1699)   
              else if (local_pf_num==0 && local_vf_num ==1700 && local_vf_active==1) `toggle_tready(1700)   
              else if (local_pf_num==0 && local_vf_num ==1701 && local_vf_active==1) `toggle_tready(1701)   
              else if (local_pf_num==0 && local_vf_num ==1702 && local_vf_active==1) `toggle_tready(1702)   
              else if (local_pf_num==0 && local_vf_num ==1703 && local_vf_active==1) `toggle_tready(1703)   
              else if (local_pf_num==0 && local_vf_num ==1704 && local_vf_active==1) `toggle_tready(1704)   
              else if (local_pf_num==0 && local_vf_num ==1705 && local_vf_active==1) `toggle_tready(1705)   
              else if (local_pf_num==0 && local_vf_num ==1706 && local_vf_active==1) `toggle_tready(1706)   
              else if (local_pf_num==0 && local_vf_num ==1707 && local_vf_active==1) `toggle_tready(1707)   
              else if (local_pf_num==0 && local_vf_num ==1708 && local_vf_active==1) `toggle_tready(1708)   
              else if (local_pf_num==0 && local_vf_num ==1709 && local_vf_active==1) `toggle_tready(1709)   
              else if (local_pf_num==0 && local_vf_num ==1710 && local_vf_active==1) `toggle_tready(1710)   
              else if (local_pf_num==0 && local_vf_num ==1711 && local_vf_active==1) `toggle_tready(1711)   
              else if (local_pf_num==0 && local_vf_num ==1712 && local_vf_active==1) `toggle_tready(1712)   
              else if (local_pf_num==0 && local_vf_num ==1713 && local_vf_active==1) `toggle_tready(1713)   
              else if (local_pf_num==0 && local_vf_num ==1714 && local_vf_active==1) `toggle_tready(1714)   
              else if (local_pf_num==0 && local_vf_num ==1715 && local_vf_active==1) `toggle_tready(1715)   
              else if (local_pf_num==0 && local_vf_num ==1716 && local_vf_active==1) `toggle_tready(1716)   
              else if (local_pf_num==0 && local_vf_num ==1717 && local_vf_active==1) `toggle_tready(1717)   
              else if (local_pf_num==0 && local_vf_num ==1718 && local_vf_active==1) `toggle_tready(1718)   
              else if (local_pf_num==0 && local_vf_num ==1719 && local_vf_active==1) `toggle_tready(1719)   
              else if (local_pf_num==0 && local_vf_num ==1720 && local_vf_active==1) `toggle_tready(1720)   
              else if (local_pf_num==0 && local_vf_num ==1721 && local_vf_active==1) `toggle_tready(1721)   
              else if (local_pf_num==0 && local_vf_num ==1722 && local_vf_active==1) `toggle_tready(1722)   
              else if (local_pf_num==0 && local_vf_num ==1723 && local_vf_active==1) `toggle_tready(1723)   
              else if (local_pf_num==0 && local_vf_num ==1724 && local_vf_active==1) `toggle_tready(1724)   
              else if (local_pf_num==0 && local_vf_num ==1725 && local_vf_active==1) `toggle_tready(1725)   
              else if (local_pf_num==0 && local_vf_num ==1726 && local_vf_active==1) `toggle_tready(1726)   
              else if (local_pf_num==0 && local_vf_num ==1727 && local_vf_active==1) `toggle_tready(1727)   
              else if (local_pf_num==0 && local_vf_num ==1728 && local_vf_active==1) `toggle_tready(1728)   
              else if (local_pf_num==0 && local_vf_num ==1729 && local_vf_active==1) `toggle_tready(1729)   
              else if (local_pf_num==0 && local_vf_num ==1730 && local_vf_active==1) `toggle_tready(1730)   
              else if (local_pf_num==0 && local_vf_num ==1731 && local_vf_active==1) `toggle_tready(1731)   
              else if (local_pf_num==0 && local_vf_num ==1732 && local_vf_active==1) `toggle_tready(1732)   
              else if (local_pf_num==0 && local_vf_num ==1733 && local_vf_active==1) `toggle_tready(1733)   
              else if (local_pf_num==0 && local_vf_num ==1734 && local_vf_active==1) `toggle_tready(1734)   
              else if (local_pf_num==0 && local_vf_num ==1735 && local_vf_active==1) `toggle_tready(1735)   
              else if (local_pf_num==0 && local_vf_num ==1736 && local_vf_active==1) `toggle_tready(1736)   
              else if (local_pf_num==0 && local_vf_num ==1737 && local_vf_active==1) `toggle_tready(1737)   
              else if (local_pf_num==0 && local_vf_num ==1738 && local_vf_active==1) `toggle_tready(1738)   
              else if (local_pf_num==0 && local_vf_num ==1739 && local_vf_active==1) `toggle_tready(1739)   
              else if (local_pf_num==0 && local_vf_num ==1740 && local_vf_active==1) `toggle_tready(1740)   
              else if (local_pf_num==0 && local_vf_num ==1741 && local_vf_active==1) `toggle_tready(1741)   
              else if (local_pf_num==0 && local_vf_num ==1742 && local_vf_active==1) `toggle_tready(1742)   
              else if (local_pf_num==0 && local_vf_num ==1743 && local_vf_active==1) `toggle_tready(1743)   
              else if (local_pf_num==0 && local_vf_num ==1744 && local_vf_active==1) `toggle_tready(1744)   
              else if (local_pf_num==0 && local_vf_num ==1745 && local_vf_active==1) `toggle_tready(1745)   
              else if (local_pf_num==0 && local_vf_num ==1746 && local_vf_active==1) `toggle_tready(1746)   
              else if (local_pf_num==0 && local_vf_num ==1747 && local_vf_active==1) `toggle_tready(1747)   
              else if (local_pf_num==0 && local_vf_num ==1748 && local_vf_active==1) `toggle_tready(1748)   
              else if (local_pf_num==0 && local_vf_num ==1749 && local_vf_active==1) `toggle_tready(1749)   
              else if (local_pf_num==0 && local_vf_num ==1750 && local_vf_active==1) `toggle_tready(1750)   
              else if (local_pf_num==0 && local_vf_num ==1751 && local_vf_active==1) `toggle_tready(1751)   
              else if (local_pf_num==0 && local_vf_num ==1752 && local_vf_active==1) `toggle_tready(1752)   
              else if (local_pf_num==0 && local_vf_num ==1753 && local_vf_active==1) `toggle_tready(1753)   
              else if (local_pf_num==0 && local_vf_num ==1754 && local_vf_active==1) `toggle_tready(1754)   
              else if (local_pf_num==0 && local_vf_num ==1755 && local_vf_active==1) `toggle_tready(1755)   
              else if (local_pf_num==0 && local_vf_num ==1756 && local_vf_active==1) `toggle_tready(1756)   
              else if (local_pf_num==0 && local_vf_num ==1757 && local_vf_active==1) `toggle_tready(1757)   
              else if (local_pf_num==0 && local_vf_num ==1758 && local_vf_active==1) `toggle_tready(1758)   
              else if (local_pf_num==0 && local_vf_num ==1759 && local_vf_active==1) `toggle_tready(1759)   
              else if (local_pf_num==0 && local_vf_num ==1760 && local_vf_active==1) `toggle_tready(1760)   
              else if (local_pf_num==0 && local_vf_num ==1761 && local_vf_active==1) `toggle_tready(1761)   
              else if (local_pf_num==0 && local_vf_num ==1762 && local_vf_active==1) `toggle_tready(1762)   
              else if (local_pf_num==0 && local_vf_num ==1763 && local_vf_active==1) `toggle_tready(1763)   
              else if (local_pf_num==0 && local_vf_num ==1764 && local_vf_active==1) `toggle_tready(1764)   
              else if (local_pf_num==0 && local_vf_num ==1765 && local_vf_active==1) `toggle_tready(1765)   
              else if (local_pf_num==0 && local_vf_num ==1766 && local_vf_active==1) `toggle_tready(1766)   
              else if (local_pf_num==0 && local_vf_num ==1767 && local_vf_active==1) `toggle_tready(1767)   
              else if (local_pf_num==0 && local_vf_num ==1768 && local_vf_active==1) `toggle_tready(1768)   
              else if (local_pf_num==0 && local_vf_num ==1769 && local_vf_active==1) `toggle_tready(1769)   
              else if (local_pf_num==0 && local_vf_num ==1770 && local_vf_active==1) `toggle_tready(1770)   
              else if (local_pf_num==0 && local_vf_num ==1771 && local_vf_active==1) `toggle_tready(1771)   
              else if (local_pf_num==0 && local_vf_num ==1772 && local_vf_active==1) `toggle_tready(1772)   
              else if (local_pf_num==0 && local_vf_num ==1773 && local_vf_active==1) `toggle_tready(1773)   
              else if (local_pf_num==0 && local_vf_num ==1774 && local_vf_active==1) `toggle_tready(1774)   
              else if (local_pf_num==0 && local_vf_num ==1775 && local_vf_active==1) `toggle_tready(1775)   
              else if (local_pf_num==0 && local_vf_num ==1776 && local_vf_active==1) `toggle_tready(1776)   
              else if (local_pf_num==0 && local_vf_num ==1777 && local_vf_active==1) `toggle_tready(1777)   
              else if (local_pf_num==0 && local_vf_num ==1778 && local_vf_active==1) `toggle_tready(1778)   
              else if (local_pf_num==0 && local_vf_num ==1779 && local_vf_active==1) `toggle_tready(1779)   
              else if (local_pf_num==0 && local_vf_num ==1780 && local_vf_active==1) `toggle_tready(1780)   
              else if (local_pf_num==0 && local_vf_num ==1781 && local_vf_active==1) `toggle_tready(1781)   
              else if (local_pf_num==0 && local_vf_num ==1782 && local_vf_active==1) `toggle_tready(1782)   
              else if (local_pf_num==0 && local_vf_num ==1783 && local_vf_active==1) `toggle_tready(1783)   
              else if (local_pf_num==0 && local_vf_num ==1784 && local_vf_active==1) `toggle_tready(1784)   
              else if (local_pf_num==0 && local_vf_num ==1785 && local_vf_active==1) `toggle_tready(1785)   
              else if (local_pf_num==0 && local_vf_num ==1786 && local_vf_active==1) `toggle_tready(1786)   
              else if (local_pf_num==0 && local_vf_num ==1787 && local_vf_active==1) `toggle_tready(1787)   
              else if (local_pf_num==0 && local_vf_num ==1788 && local_vf_active==1) `toggle_tready(1788)   
              else if (local_pf_num==0 && local_vf_num ==1789 && local_vf_active==1) `toggle_tready(1789)   
              else if (local_pf_num==0 && local_vf_num ==1790 && local_vf_active==1) `toggle_tready(1790)   
              else if (local_pf_num==0 && local_vf_num ==1791 && local_vf_active==1) `toggle_tready(1791)   
              else if (local_pf_num==0 && local_vf_num ==1792 && local_vf_active==1) `toggle_tready(1792)   
              else if (local_pf_num==0 && local_vf_num ==1793 && local_vf_active==1) `toggle_tready(1793)   
              else if (local_pf_num==0 && local_vf_num ==1794 && local_vf_active==1) `toggle_tready(1794)   
              else if (local_pf_num==0 && local_vf_num ==1795 && local_vf_active==1) `toggle_tready(1795)   
              else if (local_pf_num==0 && local_vf_num ==1796 && local_vf_active==1) `toggle_tready(1796)   
              else if (local_pf_num==0 && local_vf_num ==1797 && local_vf_active==1) `toggle_tready(1797)   
              else if (local_pf_num==0 && local_vf_num ==1798 && local_vf_active==1) `toggle_tready(1798)   
              else if (local_pf_num==0 && local_vf_num ==1799 && local_vf_active==1) `toggle_tready(1799)   
              else if (local_pf_num==0 && local_vf_num ==1800 && local_vf_active==1) `toggle_tready(1800)   
              else if (local_pf_num==0 && local_vf_num ==1801 && local_vf_active==1) `toggle_tready(1801)   
              else if (local_pf_num==0 && local_vf_num ==1802 && local_vf_active==1) `toggle_tready(1802)   
              else if (local_pf_num==0 && local_vf_num ==1803 && local_vf_active==1) `toggle_tready(1803)   
              else if (local_pf_num==0 && local_vf_num ==1804 && local_vf_active==1) `toggle_tready(1804)   
              else if (local_pf_num==0 && local_vf_num ==1805 && local_vf_active==1) `toggle_tready(1805)   
              else if (local_pf_num==0 && local_vf_num ==1806 && local_vf_active==1) `toggle_tready(1806)   
              else if (local_pf_num==0 && local_vf_num ==1807 && local_vf_active==1) `toggle_tready(1807)   
              else if (local_pf_num==0 && local_vf_num ==1808 && local_vf_active==1) `toggle_tready(1808)   
              else if (local_pf_num==0 && local_vf_num ==1809 && local_vf_active==1) `toggle_tready(1809)   
              else if (local_pf_num==0 && local_vf_num ==1810 && local_vf_active==1) `toggle_tready(1810)   
              else if (local_pf_num==0 && local_vf_num ==1811 && local_vf_active==1) `toggle_tready(1811)   
              else if (local_pf_num==0 && local_vf_num ==1812 && local_vf_active==1) `toggle_tready(1812)   
              else if (local_pf_num==0 && local_vf_num ==1813 && local_vf_active==1) `toggle_tready(1813)   
              else if (local_pf_num==0 && local_vf_num ==1814 && local_vf_active==1) `toggle_tready(1814)   
              else if (local_pf_num==0 && local_vf_num ==1815 && local_vf_active==1) `toggle_tready(1815)   
              else if (local_pf_num==0 && local_vf_num ==1816 && local_vf_active==1) `toggle_tready(1816)   
              else if (local_pf_num==0 && local_vf_num ==1817 && local_vf_active==1) `toggle_tready(1817)   
              else if (local_pf_num==0 && local_vf_num ==1818 && local_vf_active==1) `toggle_tready(1818)   
              else if (local_pf_num==0 && local_vf_num ==1819 && local_vf_active==1) `toggle_tready(1819)   
              else if (local_pf_num==0 && local_vf_num ==1820 && local_vf_active==1) `toggle_tready(1820)   
              else if (local_pf_num==0 && local_vf_num ==1821 && local_vf_active==1) `toggle_tready(1821)   
              else if (local_pf_num==0 && local_vf_num ==1822 && local_vf_active==1) `toggle_tready(1822)   
              else if (local_pf_num==0 && local_vf_num ==1823 && local_vf_active==1) `toggle_tready(1823)   
              else if (local_pf_num==0 && local_vf_num ==1824 && local_vf_active==1) `toggle_tready(1824)   
              else if (local_pf_num==0 && local_vf_num ==1825 && local_vf_active==1) `toggle_tready(1825)   
              else if (local_pf_num==0 && local_vf_num ==1826 && local_vf_active==1) `toggle_tready(1826)   
              else if (local_pf_num==0 && local_vf_num ==1827 && local_vf_active==1) `toggle_tready(1827)   
              else if (local_pf_num==0 && local_vf_num ==1828 && local_vf_active==1) `toggle_tready(1828)   
              else if (local_pf_num==0 && local_vf_num ==1829 && local_vf_active==1) `toggle_tready(1829)   
              else if (local_pf_num==0 && local_vf_num ==1830 && local_vf_active==1) `toggle_tready(1830)   
              else if (local_pf_num==0 && local_vf_num ==1831 && local_vf_active==1) `toggle_tready(1831)   
              else if (local_pf_num==0 && local_vf_num ==1832 && local_vf_active==1) `toggle_tready(1832)   
              else if (local_pf_num==0 && local_vf_num ==1833 && local_vf_active==1) `toggle_tready(1833)   
              else if (local_pf_num==0 && local_vf_num ==1834 && local_vf_active==1) `toggle_tready(1834)   
              else if (local_pf_num==0 && local_vf_num ==1835 && local_vf_active==1) `toggle_tready(1835)   
              else if (local_pf_num==0 && local_vf_num ==1836 && local_vf_active==1) `toggle_tready(1836)   
              else if (local_pf_num==0 && local_vf_num ==1837 && local_vf_active==1) `toggle_tready(1837)   
              else if (local_pf_num==0 && local_vf_num ==1838 && local_vf_active==1) `toggle_tready(1838)   
              else if (local_pf_num==0 && local_vf_num ==1839 && local_vf_active==1) `toggle_tready(1839)   
              else if (local_pf_num==0 && local_vf_num ==1840 && local_vf_active==1) `toggle_tready(1840)   
              else if (local_pf_num==0 && local_vf_num ==1841 && local_vf_active==1) `toggle_tready(1841)   
              else if (local_pf_num==0 && local_vf_num ==1842 && local_vf_active==1) `toggle_tready(1842)   
              else if (local_pf_num==0 && local_vf_num ==1843 && local_vf_active==1) `toggle_tready(1843)   
              else if (local_pf_num==0 && local_vf_num ==1844 && local_vf_active==1) `toggle_tready(1844)   
              else if (local_pf_num==0 && local_vf_num ==1845 && local_vf_active==1) `toggle_tready(1845)   
              else if (local_pf_num==0 && local_vf_num ==1846 && local_vf_active==1) `toggle_tready(1846)   
              else if (local_pf_num==0 && local_vf_num ==1847 && local_vf_active==1) `toggle_tready(1847)   
              else if (local_pf_num==0 && local_vf_num ==1848 && local_vf_active==1) `toggle_tready(1848)   
              else if (local_pf_num==0 && local_vf_num ==1849 && local_vf_active==1) `toggle_tready(1849)   
              else if (local_pf_num==0 && local_vf_num ==1850 && local_vf_active==1) `toggle_tready(1850)   
              else if (local_pf_num==0 && local_vf_num ==1851 && local_vf_active==1) `toggle_tready(1851)   
              else if (local_pf_num==0 && local_vf_num ==1852 && local_vf_active==1) `toggle_tready(1852)   
              else if (local_pf_num==0 && local_vf_num ==1853 && local_vf_active==1) `toggle_tready(1853)   
              else if (local_pf_num==0 && local_vf_num ==1854 && local_vf_active==1) `toggle_tready(1854)   
              else if (local_pf_num==0 && local_vf_num ==1855 && local_vf_active==1) `toggle_tready(1855)   
              else if (local_pf_num==0 && local_vf_num ==1856 && local_vf_active==1) `toggle_tready(1856)   
              else if (local_pf_num==0 && local_vf_num ==1857 && local_vf_active==1) `toggle_tready(1857)   
              else if (local_pf_num==0 && local_vf_num ==1858 && local_vf_active==1) `toggle_tready(1858)   
              else if (local_pf_num==0 && local_vf_num ==1859 && local_vf_active==1) `toggle_tready(1859)   
              else if (local_pf_num==0 && local_vf_num ==1860 && local_vf_active==1) `toggle_tready(1860)   
              else if (local_pf_num==0 && local_vf_num ==1861 && local_vf_active==1) `toggle_tready(1861)   
              else if (local_pf_num==0 && local_vf_num ==1862 && local_vf_active==1) `toggle_tready(1862)   
              else if (local_pf_num==0 && local_vf_num ==1863 && local_vf_active==1) `toggle_tready(1863)   
              else if (local_pf_num==0 && local_vf_num ==1864 && local_vf_active==1) `toggle_tready(1864)   
              else if (local_pf_num==0 && local_vf_num ==1865 && local_vf_active==1) `toggle_tready(1865)   
              else if (local_pf_num==0 && local_vf_num ==1866 && local_vf_active==1) `toggle_tready(1866)   
              else if (local_pf_num==0 && local_vf_num ==1867 && local_vf_active==1) `toggle_tready(1867)   
              else if (local_pf_num==0 && local_vf_num ==1868 && local_vf_active==1) `toggle_tready(1868)   
              else if (local_pf_num==0 && local_vf_num ==1869 && local_vf_active==1) `toggle_tready(1869)   
              else if (local_pf_num==0 && local_vf_num ==1870 && local_vf_active==1) `toggle_tready(1870)   
              else if (local_pf_num==0 && local_vf_num ==1871 && local_vf_active==1) `toggle_tready(1871)   
              else if (local_pf_num==0 && local_vf_num ==1872 && local_vf_active==1) `toggle_tready(1872)   
              else if (local_pf_num==0 && local_vf_num ==1873 && local_vf_active==1) `toggle_tready(1873)   
              else if (local_pf_num==0 && local_vf_num ==1874 && local_vf_active==1) `toggle_tready(1874)   
              else if (local_pf_num==0 && local_vf_num ==1875 && local_vf_active==1) `toggle_tready(1875)   
              else if (local_pf_num==0 && local_vf_num ==1876 && local_vf_active==1) `toggle_tready(1876)   
              else if (local_pf_num==0 && local_vf_num ==1877 && local_vf_active==1) `toggle_tready(1877)   
              else if (local_pf_num==0 && local_vf_num ==1878 && local_vf_active==1) `toggle_tready(1878)   
              else if (local_pf_num==0 && local_vf_num ==1879 && local_vf_active==1) `toggle_tready(1879)   
              else if (local_pf_num==0 && local_vf_num ==1880 && local_vf_active==1) `toggle_tready(1880)   
              else if (local_pf_num==0 && local_vf_num ==1881 && local_vf_active==1) `toggle_tready(1881)   
              else if (local_pf_num==0 && local_vf_num ==1882 && local_vf_active==1) `toggle_tready(1882)   
              else if (local_pf_num==0 && local_vf_num ==1883 && local_vf_active==1) `toggle_tready(1883)   
              else if (local_pf_num==0 && local_vf_num ==1884 && local_vf_active==1) `toggle_tready(1884)   
              else if (local_pf_num==0 && local_vf_num ==1885 && local_vf_active==1) `toggle_tready(1885)   
              else if (local_pf_num==0 && local_vf_num ==1886 && local_vf_active==1) `toggle_tready(1886)   
              else if (local_pf_num==0 && local_vf_num ==1887 && local_vf_active==1) `toggle_tready(1887)   
              else if (local_pf_num==0 && local_vf_num ==1888 && local_vf_active==1) `toggle_tready(1888)   
              else if (local_pf_num==0 && local_vf_num ==1889 && local_vf_active==1) `toggle_tready(1889)   
              else if (local_pf_num==0 && local_vf_num ==1890 && local_vf_active==1) `toggle_tready(1890)   
              else if (local_pf_num==0 && local_vf_num ==1891 && local_vf_active==1) `toggle_tready(1891)   
              else if (local_pf_num==0 && local_vf_num ==1892 && local_vf_active==1) `toggle_tready(1892)   
              else if (local_pf_num==0 && local_vf_num ==1893 && local_vf_active==1) `toggle_tready(1893)   
              else if (local_pf_num==0 && local_vf_num ==1894 && local_vf_active==1) `toggle_tready(1894)   
              else if (local_pf_num==0 && local_vf_num ==1895 && local_vf_active==1) `toggle_tready(1895)   
              else if (local_pf_num==0 && local_vf_num ==1896 && local_vf_active==1) `toggle_tready(1896)   
              else if (local_pf_num==0 && local_vf_num ==1897 && local_vf_active==1) `toggle_tready(1897)   
              else if (local_pf_num==0 && local_vf_num ==1898 && local_vf_active==1) `toggle_tready(1898)   
              else if (local_pf_num==0 && local_vf_num ==1899 && local_vf_active==1) `toggle_tready(1899)   
              else if (local_pf_num==0 && local_vf_num ==1900 && local_vf_active==1) `toggle_tready(1900)   
              else if (local_pf_num==0 && local_vf_num ==1901 && local_vf_active==1) `toggle_tready(1901)   
              else if (local_pf_num==0 && local_vf_num ==1902 && local_vf_active==1) `toggle_tready(1902)   
              else if (local_pf_num==0 && local_vf_num ==1903 && local_vf_active==1) `toggle_tready(1903)   
              else if (local_pf_num==0 && local_vf_num ==1904 && local_vf_active==1) `toggle_tready(1904)   
              else if (local_pf_num==0 && local_vf_num ==1905 && local_vf_active==1) `toggle_tready(1905)   
              else if (local_pf_num==0 && local_vf_num ==1906 && local_vf_active==1) `toggle_tready(1906)   
              else if (local_pf_num==0 && local_vf_num ==1907 && local_vf_active==1) `toggle_tready(1907)   
              else if (local_pf_num==0 && local_vf_num ==1908 && local_vf_active==1) `toggle_tready(1908)   
              else if (local_pf_num==0 && local_vf_num ==1909 && local_vf_active==1) `toggle_tready(1909)   
              else if (local_pf_num==0 && local_vf_num ==1910 && local_vf_active==1) `toggle_tready(1910)   
              else if (local_pf_num==0 && local_vf_num ==1911 && local_vf_active==1) `toggle_tready(1911)   
              else if (local_pf_num==0 && local_vf_num ==1912 && local_vf_active==1) `toggle_tready(1912)   
              else if (local_pf_num==0 && local_vf_num ==1913 && local_vf_active==1) `toggle_tready(1913)   
              else if (local_pf_num==0 && local_vf_num ==1914 && local_vf_active==1) `toggle_tready(1914)   
              else if (local_pf_num==0 && local_vf_num ==1915 && local_vf_active==1) `toggle_tready(1915)   
              else if (local_pf_num==0 && local_vf_num ==1916 && local_vf_active==1) `toggle_tready(1916)   
              else if (local_pf_num==0 && local_vf_num ==1917 && local_vf_active==1) `toggle_tready(1917)   
              else if (local_pf_num==0 && local_vf_num ==1918 && local_vf_active==1) `toggle_tready(1918)   
              else if (local_pf_num==0 && local_vf_num ==1919 && local_vf_active==1) `toggle_tready(1919)   
              else if (local_pf_num==0 && local_vf_num ==1920 && local_vf_active==1) `toggle_tready(1920)   
              else if (local_pf_num==0 && local_vf_num ==1921 && local_vf_active==1) `toggle_tready(1921)   
              else if (local_pf_num==0 && local_vf_num ==1922 && local_vf_active==1) `toggle_tready(1922)   
              else if (local_pf_num==0 && local_vf_num ==1923 && local_vf_active==1) `toggle_tready(1923)   
              else if (local_pf_num==0 && local_vf_num ==1924 && local_vf_active==1) `toggle_tready(1924)   
              else if (local_pf_num==0 && local_vf_num ==1925 && local_vf_active==1) `toggle_tready(1925)   
              else if (local_pf_num==0 && local_vf_num ==1926 && local_vf_active==1) `toggle_tready(1926)   
              else if (local_pf_num==0 && local_vf_num ==1927 && local_vf_active==1) `toggle_tready(1927)   
              else if (local_pf_num==0 && local_vf_num ==1928 && local_vf_active==1) `toggle_tready(1928)   
              else if (local_pf_num==0 && local_vf_num ==1929 && local_vf_active==1) `toggle_tready(1929)   
              else if (local_pf_num==0 && local_vf_num ==1930 && local_vf_active==1) `toggle_tready(1930)   
              else if (local_pf_num==0 && local_vf_num ==1931 && local_vf_active==1) `toggle_tready(1931)   
              else if (local_pf_num==0 && local_vf_num ==1932 && local_vf_active==1) `toggle_tready(1932)   
              else if (local_pf_num==0 && local_vf_num ==1933 && local_vf_active==1) `toggle_tready(1933)   
              else if (local_pf_num==0 && local_vf_num ==1934 && local_vf_active==1) `toggle_tready(1934)   
              else if (local_pf_num==0 && local_vf_num ==1935 && local_vf_active==1) `toggle_tready(1935)   
              else if (local_pf_num==0 && local_vf_num ==1936 && local_vf_active==1) `toggle_tready(1936)   
              else if (local_pf_num==0 && local_vf_num ==1937 && local_vf_active==1) `toggle_tready(1937)   
              else if (local_pf_num==0 && local_vf_num ==1938 && local_vf_active==1) `toggle_tready(1938)   
              else if (local_pf_num==0 && local_vf_num ==1939 && local_vf_active==1) `toggle_tready(1939)   
              else if (local_pf_num==0 && local_vf_num ==1940 && local_vf_active==1) `toggle_tready(1940)   
              else if (local_pf_num==0 && local_vf_num ==1941 && local_vf_active==1) `toggle_tready(1941)   
              else if (local_pf_num==0 && local_vf_num ==1942 && local_vf_active==1) `toggle_tready(1942)   
              else if (local_pf_num==0 && local_vf_num ==1943 && local_vf_active==1) `toggle_tready(1943)   
              else if (local_pf_num==0 && local_vf_num ==1944 && local_vf_active==1) `toggle_tready(1944)   
              else if (local_pf_num==0 && local_vf_num ==1945 && local_vf_active==1) `toggle_tready(1945)   
              else if (local_pf_num==0 && local_vf_num ==1946 && local_vf_active==1) `toggle_tready(1946)   
              else if (local_pf_num==0 && local_vf_num ==1947 && local_vf_active==1) `toggle_tready(1947)   
              else if (local_pf_num==0 && local_vf_num ==1948 && local_vf_active==1) `toggle_tready(1948)   
              else if (local_pf_num==0 && local_vf_num ==1949 && local_vf_active==1) `toggle_tready(1949)   
              else if (local_pf_num==0 && local_vf_num ==1950 && local_vf_active==1) `toggle_tready(1950)   
              else if (local_pf_num==0 && local_vf_num ==1951 && local_vf_active==1) `toggle_tready(1951)   
              else if (local_pf_num==0 && local_vf_num ==1952 && local_vf_active==1) `toggle_tready(1952)   
              else if (local_pf_num==0 && local_vf_num ==1953 && local_vf_active==1) `toggle_tready(1953)   
              else if (local_pf_num==0 && local_vf_num ==1954 && local_vf_active==1) `toggle_tready(1954)   
              else if (local_pf_num==0 && local_vf_num ==1955 && local_vf_active==1) `toggle_tready(1955)   
              else if (local_pf_num==0 && local_vf_num ==1956 && local_vf_active==1) `toggle_tready(1956)   
              else if (local_pf_num==0 && local_vf_num ==1957 && local_vf_active==1) `toggle_tready(1957)   
              else if (local_pf_num==0 && local_vf_num ==1958 && local_vf_active==1) `toggle_tready(1958)   
              else if (local_pf_num==0 && local_vf_num ==1959 && local_vf_active==1) `toggle_tready(1959)   
              else if (local_pf_num==0 && local_vf_num ==1960 && local_vf_active==1) `toggle_tready(1960)   
              else if (local_pf_num==0 && local_vf_num ==1961 && local_vf_active==1) `toggle_tready(1961)   
              else if (local_pf_num==0 && local_vf_num ==1962 && local_vf_active==1) `toggle_tready(1962)   
              else if (local_pf_num==0 && local_vf_num ==1963 && local_vf_active==1) `toggle_tready(1963)   
              else if (local_pf_num==0 && local_vf_num ==1964 && local_vf_active==1) `toggle_tready(1964)   
              else if (local_pf_num==0 && local_vf_num ==1965 && local_vf_active==1) `toggle_tready(1965)   
              else if (local_pf_num==0 && local_vf_num ==1966 && local_vf_active==1) `toggle_tready(1966)   
              else if (local_pf_num==0 && local_vf_num ==1967 && local_vf_active==1) `toggle_tready(1967)   
              else if (local_pf_num==0 && local_vf_num ==1968 && local_vf_active==1) `toggle_tready(1968)   
              else if (local_pf_num==0 && local_vf_num ==1969 && local_vf_active==1) `toggle_tready(1969)   
              else if (local_pf_num==0 && local_vf_num ==1970 && local_vf_active==1) `toggle_tready(1970)   
              else if (local_pf_num==0 && local_vf_num ==1971 && local_vf_active==1) `toggle_tready(1971)   
              else if (local_pf_num==0 && local_vf_num ==1972 && local_vf_active==1) `toggle_tready(1972)   
              else if (local_pf_num==0 && local_vf_num ==1973 && local_vf_active==1) `toggle_tready(1973)   
              else if (local_pf_num==0 && local_vf_num ==1974 && local_vf_active==1) `toggle_tready(1974)   
              else if (local_pf_num==0 && local_vf_num ==1975 && local_vf_active==1) `toggle_tready(1975)   
              else if (local_pf_num==0 && local_vf_num ==1976 && local_vf_active==1) `toggle_tready(1976)   
              else if (local_pf_num==0 && local_vf_num ==1977 && local_vf_active==1) `toggle_tready(1977)   
              else if (local_pf_num==0 && local_vf_num ==1978 && local_vf_active==1) `toggle_tready(1978)   
              else if (local_pf_num==0 && local_vf_num ==1979 && local_vf_active==1) `toggle_tready(1979)   
              else if (local_pf_num==0 && local_vf_num ==1980 && local_vf_active==1) `toggle_tready(1980)   
              else if (local_pf_num==0 && local_vf_num ==1981 && local_vf_active==1) `toggle_tready(1981)   
              else if (local_pf_num==0 && local_vf_num ==1982 && local_vf_active==1) `toggle_tready(1982)   
              else if (local_pf_num==0 && local_vf_num ==1983 && local_vf_active==1) `toggle_tready(1983)   
              else if (local_pf_num==0 && local_vf_num ==1984 && local_vf_active==1) `toggle_tready(1984)   
              else if (local_pf_num==0 && local_vf_num ==1985 && local_vf_active==1) `toggle_tready(1985)   
              else if (local_pf_num==0 && local_vf_num ==1986 && local_vf_active==1) `toggle_tready(1986)   
              else if (local_pf_num==0 && local_vf_num ==1987 && local_vf_active==1) `toggle_tready(1987)   
              else if (local_pf_num==0 && local_vf_num ==1988 && local_vf_active==1) `toggle_tready(1988)   
              else if (local_pf_num==0 && local_vf_num ==1989 && local_vf_active==1) `toggle_tready(1989)   
              else if (local_pf_num==0 && local_vf_num ==1990 && local_vf_active==1) `toggle_tready(1990)   
              else if (local_pf_num==0 && local_vf_num ==1991 && local_vf_active==1) `toggle_tready(1991)   
              else if (local_pf_num==0 && local_vf_num ==1992 && local_vf_active==1) `toggle_tready(1992)   
              else if (local_pf_num==0 && local_vf_num ==1993 && local_vf_active==1) `toggle_tready(1993)   
              else if (local_pf_num==0 && local_vf_num ==1994 && local_vf_active==1) `toggle_tready(1994)   
              else if (local_pf_num==0 && local_vf_num ==1995 && local_vf_active==1) `toggle_tready(1995)   
              else if (local_pf_num==0 && local_vf_num ==1996 && local_vf_active==1) `toggle_tready(1996)   
              else if (local_pf_num==0 && local_vf_num ==1997 && local_vf_active==1) `toggle_tready(1997)   
              else if (local_pf_num==0 && local_vf_num ==1998 && local_vf_active==1) `toggle_tready(1998)   
              else if (local_pf_num==0 && local_vf_num ==1999 && local_vf_active==1) `toggle_tready(1999)   
              else if (local_pf_num==0 && local_vf_num ==2000 && local_vf_active==1) `toggle_tready(2000)   
              else if (local_pf_num==0 && local_vf_num ==2001 && local_vf_active==1) `toggle_tready(2001)   
              else if (local_pf_num==0 && local_vf_num ==2002 && local_vf_active==1) `toggle_tready(2002)   
              else if (local_pf_num==0 && local_vf_num ==2003 && local_vf_active==1) `toggle_tready(2003)   
              else if (local_pf_num==0 && local_vf_num ==2004 && local_vf_active==1) `toggle_tready(2004)   
              else if (local_pf_num==0 && local_vf_num ==2005 && local_vf_active==1) `toggle_tready(2005)   
              else if (local_pf_num==0 && local_vf_num ==2006 && local_vf_active==1) `toggle_tready(2006)   
              else if (local_pf_num==0 && local_vf_num ==2007 && local_vf_active==1) `toggle_tready(2007)   
              else if (local_pf_num==0 && local_vf_num ==2008 && local_vf_active==1) `toggle_tready(2008)   
              else if (local_pf_num==0 && local_vf_num ==2009 && local_vf_active==1) `toggle_tready(2009)   
              else if (local_pf_num==0 && local_vf_num ==2010 && local_vf_active==1) `toggle_tready(2010)   
              else if (local_pf_num==0 && local_vf_num ==2011 && local_vf_active==1) `toggle_tready(2011)   
              else if (local_pf_num==0 && local_vf_num ==2012 && local_vf_active==1) `toggle_tready(2012)   
              else if (local_pf_num==0 && local_vf_num ==2013 && local_vf_active==1) `toggle_tready(2013)   
              else if (local_pf_num==0 && local_vf_num ==2014 && local_vf_active==1) `toggle_tready(2014)   
              else if (local_pf_num==0 && local_vf_num ==2015 && local_vf_active==1) `toggle_tready(2015)   
              else if (local_pf_num==0 && local_vf_num ==2016 && local_vf_active==1) `toggle_tready(2016)   
              else if (local_pf_num==0 && local_vf_num ==2017 && local_vf_active==1) `toggle_tready(2017)   
              else if (local_pf_num==0 && local_vf_num ==2018 && local_vf_active==1) `toggle_tready(2018)   
              else if (local_pf_num==0 && local_vf_num ==2019 && local_vf_active==1) `toggle_tready(2019)   
              else if (local_pf_num==0 && local_vf_num ==2020 && local_vf_active==1) `toggle_tready(2020)   
              else if (local_pf_num==0 && local_vf_num ==2021 && local_vf_active==1) `toggle_tready(2021)   
              else if (local_pf_num==0 && local_vf_num ==2022 && local_vf_active==1) `toggle_tready(2022)   
              else if (local_pf_num==0 && local_vf_num ==2023 && local_vf_active==1) `toggle_tready(2023)   
              else if (local_pf_num==0 && local_vf_num ==2024 && local_vf_active==1) `toggle_tready(2024)   
              else if (local_pf_num==0 && local_vf_num ==2025 && local_vf_active==1) `toggle_tready(2025)   
              else if (local_pf_num==0 && local_vf_num ==2026 && local_vf_active==1) `toggle_tready(2026)   
              else if (local_pf_num==0 && local_vf_num ==2027 && local_vf_active==1) `toggle_tready(2027)   
              else if (local_pf_num==0 && local_vf_num ==2028 && local_vf_active==1) `toggle_tready(2028)   
              else if (local_pf_num==0 && local_vf_num ==2029 && local_vf_active==1) `toggle_tready(2029)   
              else if (local_pf_num==0 && local_vf_num ==2030 && local_vf_active==1) `toggle_tready(2030)   
              else if (local_pf_num==0 && local_vf_num ==2031 && local_vf_active==1) `toggle_tready(2031)   
              else if (local_pf_num==0 && local_vf_num ==2032 && local_vf_active==1) `toggle_tready(2032)   
              else if (local_pf_num==0 && local_vf_num ==2033 && local_vf_active==1) `toggle_tready(2033)   
              else if (local_pf_num==0 && local_vf_num ==2034 && local_vf_active==1) `toggle_tready(2034)   
              else if (local_pf_num==0 && local_vf_num ==2035 && local_vf_active==1) `toggle_tready(2035)   
              else if (local_pf_num==0 && local_vf_num ==2036 && local_vf_active==1) `toggle_tready(2036)   
              else if (local_pf_num==0 && local_vf_num ==2037 && local_vf_active==1) `toggle_tready(2037)   
              else if (local_pf_num==0 && local_vf_num ==2038 && local_vf_active==1) `toggle_tready(2038)   
              else if (local_pf_num==0 && local_vf_num ==2039 && local_vf_active==1) `toggle_tready(2039)   
              else if (local_pf_num==0 && local_vf_num ==2040 && local_vf_active==1) `toggle_tready(2040)   
              else if (local_pf_num==0 && local_vf_num ==2041 && local_vf_active==1) `toggle_tready(2041)   
              else if (local_pf_num==0 && local_vf_num ==2042 && local_vf_active==1) `toggle_tready(2042)   
              else if (local_pf_num==0 && local_vf_num ==2043 && local_vf_active==1) `toggle_tready(2043)   
              else if (local_pf_num==0 && local_vf_num ==2044 && local_vf_active==1) `toggle_tready(2044)   
              else if (local_pf_num==0 && local_vf_num ==2045 && local_vf_active==1) `toggle_tready(2045)   
              else if (local_pf_num==0 && local_vf_num ==2046 && local_vf_active==1) `toggle_tready(2046)   
              else if (local_pf_num==0 && local_vf_num ==2047 && local_vf_active==1) `toggle_tready(2047)   
              `endif
          end
          
            //=============================================
            // Starting request sequence on Host master
            //=============================================        
               begin
                `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_H, {tlp_length  == local_tlp_length  ;
                                                                             pf_num      == local_pf_num      ;
                                                                             vf_num      == local_vf_num      ;
                                                                             vf_active   == local_vf_active   ;
                                                                             payload     == local_payload     ;
                                                                             direction   == 1'b0              ;
                                                              })
        
               end
             join
           end
           count = 0; 
         end    
         end
      `uvm_info(get_name(), "Exiting sequence...", UVM_LOW)
    endtask : body

endclass
          
