// Copyright 2021 Intel Corporation
// SPDX-License-Identifier: MIT

`include "gram_sdp.v"
`include "ram_1r1w.sv"
`include "bfifo.sv"
`include "pfa_master.sv"
`include "pfa_master_tb.sv"
